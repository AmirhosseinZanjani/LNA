magic
tech sky130A
magscale 1 2
timestamp 1710869846
<< viali >>
rect 1117 2317 1169 2369
rect 23755 2316 23807 2368
rect -18 2102 34 2154
rect 24887 2101 24939 2153
rect -18 178 34 230
rect 24890 178 24942 230
rect 85 -17 137 35
rect 1117 -17 1169 35
rect 23755 -18 23807 34
rect 24782 -16 24834 36
<< metal1 >>
rect 1105 2369 1181 2375
rect 1105 2317 1117 2369
rect 1169 2317 1181 2369
rect 1105 2311 1181 2317
rect 23743 2368 23819 2374
rect 23743 2316 23755 2368
rect 23807 2316 23819 2368
rect 23743 2310 23819 2316
rect 1107 2213 1117 2265
rect 1169 2213 1179 2265
rect 3165 2213 3175 2265
rect 3227 2213 3237 2265
rect 5223 2213 5233 2265
rect 5285 2213 5295 2265
rect 7281 2211 7291 2263
rect 7343 2211 7353 2263
rect 9339 2213 9349 2265
rect 9401 2213 9411 2265
rect 11396 2213 11406 2265
rect 11458 2213 11468 2265
rect 13455 2213 13465 2265
rect 13517 2213 13527 2265
rect 15513 2213 15523 2265
rect 15575 2213 15585 2265
rect 17571 2213 17581 2265
rect 17633 2213 17643 2265
rect 19629 2213 19639 2265
rect 19691 2213 19701 2265
rect 21687 2213 21697 2265
rect 21749 2213 21759 2265
rect 23745 2213 23755 2265
rect 23807 2213 23817 2265
rect -30 2154 46 2160
rect -30 2102 -18 2154
rect 34 2102 46 2154
rect 75 2102 85 2154
rect 137 2102 147 2154
rect 2133 2102 2143 2154
rect 2195 2102 2205 2154
rect 4192 2102 4202 2154
rect 4254 2102 4264 2154
rect 6251 2102 6261 2154
rect 6313 2102 6323 2154
rect 8309 2102 8319 2154
rect 8371 2102 8381 2154
rect 10366 2102 10376 2154
rect 10428 2102 10438 2154
rect 12424 2102 12434 2154
rect 12486 2102 12496 2154
rect 14477 2102 14487 2154
rect 14539 2102 14549 2154
rect 16543 2102 16553 2154
rect 16605 2102 16615 2154
rect 18599 2102 18609 2154
rect 18661 2102 18671 2154
rect -30 2096 46 2102
rect 20656 2101 20666 2153
rect 20718 2101 20728 2153
rect 22717 2102 22727 2154
rect 22779 2102 22789 2154
rect 24875 2153 24951 2159
rect 24771 2101 24781 2153
rect 24833 2101 24843 2153
rect 24875 2101 24887 2153
rect 24939 2101 24951 2153
rect 24875 2095 24951 2101
rect -30 230 46 236
rect 24878 230 24954 236
rect -30 178 -18 230
rect 34 178 46 230
rect 75 178 85 230
rect 137 178 147 230
rect -30 172 46 178
rect 2133 177 2143 229
rect 2195 177 2205 229
rect 4192 177 4202 229
rect 4254 177 4264 229
rect 6250 178 6260 230
rect 6312 178 6322 230
rect 8308 178 8318 230
rect 8370 178 8380 230
rect 10366 177 10376 229
rect 10428 177 10438 229
rect 12424 177 12434 229
rect 12486 177 12496 229
rect 14478 176 14488 228
rect 14540 176 14550 228
rect 16543 176 16553 228
rect 16605 176 16615 228
rect 18601 178 18611 230
rect 18663 178 18673 230
rect 20657 178 20667 230
rect 20719 178 20729 230
rect 22716 178 22726 230
rect 22778 178 22788 230
rect 24772 178 24782 230
rect 24834 178 24844 230
rect 24878 178 24890 230
rect 24942 178 24954 230
rect 24878 172 24954 178
rect 1107 85 1117 137
rect 1169 85 1179 137
rect 3165 85 3175 137
rect 3227 85 3237 137
rect 5223 85 5233 137
rect 5285 85 5295 137
rect 7281 85 7291 137
rect 7343 85 7353 137
rect 9339 85 9349 137
rect 9401 85 9411 137
rect 11397 85 11407 137
rect 11459 85 11469 137
rect 13455 85 13465 137
rect 13517 85 13527 137
rect 15513 85 15523 137
rect 15575 85 15585 137
rect 17571 85 17581 137
rect 17633 85 17643 137
rect 19629 85 19639 137
rect 19691 85 19701 137
rect 21687 85 21697 137
rect 21749 85 21759 137
rect 23745 85 23755 137
rect 23807 85 23817 137
rect 73 35 149 41
rect 73 -17 85 35
rect 137 -17 149 35
rect 73 -23 149 -17
rect 1105 35 1181 41
rect 1105 -17 1117 35
rect 1169 -17 1181 35
rect 1105 -23 1181 -17
rect 23743 34 23819 40
rect 23743 -18 23755 34
rect 23807 -18 23819 34
rect 23743 -24 23819 -18
rect 24770 36 24846 42
rect 24770 -16 24782 36
rect 24834 -16 24846 36
rect 24770 -22 24846 -16
<< via1 >>
rect 1117 2317 1169 2369
rect 23755 2316 23807 2368
rect 1117 2213 1169 2265
rect 3175 2213 3227 2265
rect 5233 2213 5285 2265
rect 7291 2211 7343 2263
rect 9349 2213 9401 2265
rect 11406 2213 11458 2265
rect 13465 2213 13517 2265
rect 15523 2213 15575 2265
rect 17581 2213 17633 2265
rect 19639 2213 19691 2265
rect 21697 2213 21749 2265
rect 23755 2213 23807 2265
rect -18 2102 34 2154
rect 85 2102 137 2154
rect 2143 2102 2195 2154
rect 4202 2102 4254 2154
rect 6261 2102 6313 2154
rect 8319 2102 8371 2154
rect 10376 2102 10428 2154
rect 12434 2102 12486 2154
rect 14487 2102 14539 2154
rect 16553 2102 16605 2154
rect 18609 2102 18661 2154
rect 20666 2101 20718 2153
rect 22727 2102 22779 2154
rect 24781 2101 24833 2153
rect 24887 2101 24939 2153
rect -18 178 34 230
rect 85 178 137 230
rect 2143 177 2195 229
rect 4202 177 4254 229
rect 6260 178 6312 230
rect 8318 178 8370 230
rect 10376 177 10428 229
rect 12434 177 12486 229
rect 14488 176 14540 228
rect 16553 176 16605 228
rect 18611 178 18663 230
rect 20667 178 20719 230
rect 22726 178 22778 230
rect 24782 178 24834 230
rect 24890 178 24942 230
rect 1117 85 1169 137
rect 3175 85 3227 137
rect 5233 85 5285 137
rect 7291 85 7343 137
rect 9349 85 9401 137
rect 11407 85 11459 137
rect 13465 85 13517 137
rect 15523 85 15575 137
rect 17581 85 17633 137
rect 19639 85 19691 137
rect 21697 85 21749 137
rect 23755 85 23807 137
rect 85 -17 137 35
rect 1117 -17 1169 35
rect 23755 -18 23807 34
rect 24782 -16 24834 36
<< metal2 >>
rect 1117 2369 1169 3024
rect 3175 2517 3227 3024
rect 5233 2517 5285 3024
rect 7291 2517 7343 3024
rect 9349 2517 9401 3024
rect 11407 2517 11460 3024
rect 13465 2767 13517 3024
rect 13463 2757 13519 2767
rect 15523 2764 15575 3024
rect 17581 2765 17633 3024
rect 19639 2766 19691 3024
rect 13463 2691 13519 2701
rect 15520 2754 15576 2764
rect 3173 2507 3229 2517
rect 3173 2441 3229 2451
rect 5231 2507 5287 2517
rect 5231 2441 5287 2451
rect 7289 2507 7345 2517
rect 7289 2441 7345 2451
rect 9347 2507 9403 2517
rect 9347 2441 9403 2451
rect 11405 2507 11461 2517
rect 11405 2441 11461 2451
rect 1117 2265 1169 2317
rect -17 2164 137 2170
rect -18 2154 137 2164
rect 34 2102 85 2154
rect -18 2092 34 2102
rect -18 231 34 240
rect 85 231 137 2102
rect -18 230 137 231
rect 34 178 85 230
rect -18 168 137 178
rect -17 163 137 168
rect 85 35 137 163
rect 85 -553 137 -17
rect 1117 137 1169 2213
rect 3175 2265 3227 2441
rect 2143 2154 2195 2170
rect 2143 229 2195 2102
rect 1117 35 1169 85
rect 1117 -27 1169 -17
rect 2142 177 2143 179
rect 2142 67 2195 177
rect 3175 137 3227 2213
rect 5233 2265 5285 2441
rect 3175 75 3227 85
rect 4202 2154 4254 2170
rect 4202 229 4254 2102
rect 2142 -108 2194 67
rect 2140 -118 2196 -108
rect 2140 -184 2196 -174
rect 2142 -559 2194 -184
rect 4202 -234 4254 177
rect 5233 137 5285 2213
rect 7291 2263 7343 2441
rect 6261 2154 6313 2171
rect 6261 240 6313 2102
rect 6260 230 6313 240
rect 6312 178 6313 230
rect 6260 168 6313 178
rect 5233 75 5285 85
rect 6261 165 6313 168
rect 6261 67 6315 165
rect 7291 137 7343 2211
rect 9349 2265 9401 2441
rect 11407 2275 11460 2441
rect 8319 2154 8371 2170
rect 8319 240 8371 2102
rect 8318 230 8371 240
rect 8370 178 8371 230
rect 8318 168 8371 178
rect 7291 75 7343 85
rect 6263 -109 6315 67
rect 6260 -119 6316 -109
rect 6260 -185 6316 -175
rect 4199 -244 4255 -234
rect 4199 -310 4255 -300
rect 4202 -561 4254 -310
rect 6263 -573 6315 -185
rect 8319 -234 8371 168
rect 9349 137 9401 2213
rect 11406 2265 11460 2275
rect 13465 2265 13517 2691
rect 15520 2688 15576 2698
rect 17579 2755 17635 2765
rect 17579 2689 17635 2699
rect 19636 2756 19692 2766
rect 21697 2765 21749 3024
rect 19636 2690 19692 2700
rect 21694 2755 21750 2765
rect 11458 2213 11459 2265
rect 11406 2203 11459 2213
rect 9349 75 9401 85
rect 10376 2154 10428 2170
rect 10376 229 10428 2102
rect 10376 -110 10428 177
rect 11407 137 11459 2203
rect 12434 2154 12486 2171
rect 12434 229 12486 2102
rect 12434 133 12486 177
rect 11407 75 11459 85
rect 12433 67 12486 133
rect 13465 137 13517 2213
rect 15523 2265 15575 2688
rect 14487 2154 14539 2170
rect 14487 238 14539 2102
rect 14487 228 14540 238
rect 14487 176 14488 228
rect 14487 166 14540 176
rect 14487 131 14539 166
rect 10373 -120 10429 -110
rect 10373 -186 10429 -176
rect 8315 -244 8371 -234
rect 8315 -310 8371 -300
rect 8319 -659 8371 -310
rect 10376 -606 10428 -186
rect 12433 -233 12485 67
rect 13465 -110 13517 85
rect 14486 67 14539 131
rect 15523 137 15575 2213
rect 17581 2265 17633 2689
rect 13462 -120 13518 -110
rect 13462 -186 13518 -176
rect 12431 -243 12487 -233
rect 12431 -309 12487 -299
rect 12433 -605 12485 -309
rect 14486 -358 14538 67
rect 15523 -109 15575 85
rect 16553 2154 16605 2170
rect 16553 228 16605 2102
rect 15522 -119 15578 -109
rect 15522 -185 15578 -175
rect 14483 -368 14539 -358
rect 14483 -434 14539 -424
rect 14486 -607 14538 -434
rect 16553 -484 16605 176
rect 17581 137 17633 2213
rect 19639 2265 19691 2690
rect 21694 2689 21750 2699
rect 18610 2164 18662 2171
rect 18609 2154 18662 2164
rect 18661 2102 18662 2154
rect 18609 2092 18662 2102
rect 17581 -109 17633 85
rect 18610 240 18662 2092
rect 18610 230 18663 240
rect 18610 178 18611 230
rect 18610 168 18663 178
rect 17579 -119 17635 -109
rect 17579 -185 17635 -175
rect 18610 -360 18662 168
rect 19639 155 19691 2213
rect 21697 2265 21749 2689
rect 20667 2163 20719 2175
rect 20666 2153 20719 2163
rect 20718 2101 20719 2153
rect 20666 2091 20719 2101
rect 19637 137 19691 155
rect 19637 85 19639 137
rect 19637 -111 19691 85
rect 19635 -121 19691 -111
rect 19635 -187 19691 -177
rect 20667 230 20719 2091
rect 18607 -370 18663 -360
rect 18607 -436 18663 -426
rect 16546 -494 16605 -484
rect 16602 -550 16605 -494
rect 16546 -560 16605 -550
rect 16553 -609 16605 -560
rect 18610 -608 18662 -436
rect 20667 -484 20719 178
rect 21697 137 21749 2213
rect 23755 2368 23807 3024
rect 23755 2265 23807 2316
rect 22727 2154 22779 2181
rect 22727 240 22779 2102
rect 22726 230 22779 240
rect 22778 178 22779 230
rect 22726 168 22779 178
rect 21697 -109 21749 85
rect 21694 -119 21750 -109
rect 21694 -185 21750 -175
rect 22727 -360 22779 168
rect 23755 137 23807 2213
rect 24781 2153 24940 2184
rect 24833 2101 24887 2153
rect 24939 2101 24940 2153
rect 24781 2091 24834 2101
rect 24887 2091 24939 2101
rect 24782 230 24834 2091
rect 24890 230 24942 240
rect 24769 178 24782 230
rect 24834 178 24890 230
rect 24942 178 24943 230
rect 24769 162 24943 178
rect 23755 34 23807 85
rect 23755 -28 23807 -18
rect 24782 36 24834 162
rect 22723 -370 22779 -360
rect 22723 -436 22779 -426
rect 20665 -494 20721 -484
rect 20665 -560 20721 -550
rect 20667 -604 20719 -560
rect 22727 -598 22779 -436
rect 24782 -595 24834 -16
<< via2 >>
rect 13463 2701 13519 2757
rect 15520 2698 15576 2754
rect 3173 2451 3229 2507
rect 5231 2451 5287 2507
rect 7289 2451 7345 2507
rect 9347 2451 9403 2507
rect 11405 2451 11461 2507
rect 2140 -174 2196 -118
rect 6260 -175 6316 -119
rect 4199 -300 4255 -244
rect 17579 2699 17635 2755
rect 19636 2700 19692 2756
rect 21694 2699 21750 2755
rect 10373 -176 10429 -120
rect 8315 -300 8371 -244
rect 13462 -176 13518 -120
rect 12431 -299 12487 -243
rect 15522 -175 15578 -119
rect 14483 -424 14539 -368
rect 17579 -175 17635 -119
rect 19635 -177 19691 -121
rect 18607 -426 18663 -370
rect 16546 -550 16602 -494
rect 21694 -175 21750 -119
rect 22723 -426 22779 -370
rect 20665 -550 20721 -494
<< metal3 >>
rect 84 2882 1229 2883
rect 84 2822 24844 2882
rect 84 2757 1229 2758
rect 13453 2757 13529 2762
rect 15510 2757 15586 2759
rect 17569 2757 17645 2760
rect 19626 2757 19702 2761
rect 21684 2757 21760 2760
rect 84 2701 13463 2757
rect 13519 2756 24844 2757
rect 13519 2755 19636 2756
rect 13519 2754 17579 2755
rect 13519 2701 15520 2754
rect 84 2698 15520 2701
rect 15576 2699 17579 2754
rect 17635 2700 19636 2755
rect 19692 2755 24844 2756
rect 19692 2700 21694 2755
rect 17635 2699 21694 2700
rect 21750 2699 24844 2755
rect 15576 2698 24844 2699
rect 84 2697 24844 2698
rect 13453 2696 13529 2697
rect 15510 2693 15586 2697
rect 17569 2694 17645 2697
rect 19626 2695 19702 2697
rect 21684 2694 21760 2697
rect 84 2635 5348 2636
rect 84 2634 7408 2635
rect 84 2633 11539 2634
rect 84 2573 24844 2633
rect 3163 2511 3239 2512
rect 84 2509 3328 2511
rect 5221 2509 5297 2512
rect 7279 2509 7355 2512
rect 9337 2509 9413 2512
rect 11395 2509 11471 2512
rect 84 2507 24844 2509
rect 84 2451 3173 2507
rect 3229 2451 5231 2507
rect 5287 2451 7289 2507
rect 7345 2451 9347 2507
rect 9403 2451 11405 2507
rect 11461 2451 24844 2507
rect 84 2449 24844 2451
rect 3163 2446 3239 2449
rect 5221 2446 5297 2449
rect 7279 2446 7355 2449
rect 9337 2446 9413 2449
rect 11395 2446 11471 2449
rect 2130 -117 2206 -113
rect 6250 -117 6326 -114
rect 10363 -117 10439 -115
rect 13452 -117 13528 -115
rect 15512 -117 15588 -114
rect 17569 -117 17645 -114
rect 19625 -117 19701 -116
rect 21684 -117 21760 -114
rect 84 -118 24844 -117
rect 84 -174 2140 -118
rect 2196 -119 24844 -118
rect 2196 -174 6260 -119
rect 84 -175 6260 -174
rect 6316 -120 15522 -119
rect 6316 -175 10373 -120
rect 84 -176 10373 -175
rect 10429 -176 13462 -120
rect 13518 -175 15522 -120
rect 15578 -175 17579 -119
rect 17635 -121 21694 -119
rect 17635 -175 19635 -121
rect 13518 -176 19635 -175
rect 84 -177 19635 -176
rect 19691 -175 21694 -121
rect 21750 -175 24844 -119
rect 19691 -177 24844 -175
rect 84 -178 24844 -177
rect 2130 -179 2206 -178
rect 6250 -180 6326 -178
rect 10363 -181 10439 -178
rect 13452 -181 13528 -178
rect 15512 -180 15588 -178
rect 17569 -180 17645 -178
rect 19625 -182 19701 -178
rect 21684 -180 21760 -178
rect 4189 -242 4265 -239
rect 8305 -242 8381 -239
rect 12421 -242 12497 -238
rect 84 -243 24844 -242
rect 84 -244 12431 -243
rect 84 -300 4199 -244
rect 4255 -300 8315 -244
rect 8371 -299 12431 -244
rect 12487 -299 24844 -243
rect 8371 -300 24844 -299
rect 84 -303 24844 -300
rect 4189 -305 4265 -303
rect 8305 -305 8381 -303
rect 12421 -304 12497 -303
rect 14473 -367 14549 -363
rect 18597 -367 18673 -365
rect 22713 -367 22789 -365
rect 84 -368 24844 -367
rect 84 -424 14483 -368
rect 14539 -370 24844 -368
rect 14539 -424 18607 -370
rect 84 -426 18607 -424
rect 18663 -426 22723 -370
rect 22779 -426 24844 -370
rect 84 -428 24844 -426
rect 14473 -429 14549 -428
rect 18597 -431 18673 -428
rect 22713 -431 22789 -428
rect 16536 -492 16612 -489
rect 20655 -492 20731 -489
rect 84 -494 24844 -492
rect 84 -550 16546 -494
rect 16602 -550 20665 -494
rect 20721 -550 24844 -494
rect 84 -553 24844 -550
rect 16536 -555 16612 -553
rect 20655 -555 20731 -553
rect 79 -678 24844 -618
use core_pullup_m3_cell  core_pullup_m3_cell_0
timestamp 1710869429
transform 1 0 436529 0 1 -1962574
box -461540 1961077 -436441 1965497
use core_pullup_m3_cell  core_pullup_m3_cell_1
timestamp 1710869429
transform 1 0 486377 0 1 -1962574
box -461540 1961077 -436441 1965497
use sky130_fd_pr__pfet_01v8_X3BJMD  sky130_fd_pr__pfet_01v8_X3BJMD_0
timestamp 1710847391
transform 1 0 12462 0 1 1166
box -12515 -1219 12515 1219
<< end >>
