magic
tech sky130A
magscale 1 2
timestamp 1710254310
<< nwell >>
rect -1650 1348 -1358 1792
rect -1346 1526 -1340 1548
rect -1346 1492 -1250 1526
rect -1346 1476 -1340 1492
rect -1342 1454 -1340 1476
rect -1346 1348 -1340 1454
rect -1650 1228 -1340 1348
rect 484 1228 748 1794
rect -1650 1226 -1358 1228
<< psubdiff >>
rect -1596 2002 -1572 2098
rect -1384 2002 -1360 2098
rect 436 2002 460 2098
rect 648 2002 672 2098
rect -1598 918 -1574 1014
rect -1386 918 -1362 1014
rect 436 918 460 1014
rect 648 918 672 1014
<< nsubdiff >>
rect -1612 1596 -1374 1626
rect -1612 1406 -1580 1596
rect -1408 1406 -1374 1596
rect -1612 1380 -1374 1406
rect 446 1598 684 1626
rect 446 1408 480 1598
rect 652 1408 684 1598
rect 446 1380 684 1408
<< psubdiffcont >>
rect -1572 2002 -1384 2098
rect 460 2002 648 2098
rect -1574 918 -1386 1014
rect 460 918 648 1014
<< nsubdiffcont >>
rect -1580 1406 -1408 1596
rect 480 1408 652 1598
<< locali >>
rect -1588 2002 -1572 2098
rect -1384 2002 -1368 2098
rect 417 2070 432 2071
rect 417 2037 428 2070
rect 444 2002 460 2098
rect 648 2002 664 2098
rect -1606 1596 -1374 1612
rect -1606 1406 -1580 1596
rect -1408 1406 -1374 1596
rect 446 1598 680 1614
rect -1320 1492 -1250 1526
rect -1606 1390 -1374 1406
rect 446 1408 480 1598
rect 652 1408 680 1598
rect 446 1392 680 1408
rect -1590 918 -1574 1014
rect -1386 918 -1370 1014
rect 444 918 460 1014
rect 648 918 664 1014
<< viali >>
rect -478 1936 -444 1970
rect -1302 1798 -1268 1832
rect -1210 1798 -1176 1832
rect -1038 1800 -1004 1834
rect -946 1800 -912 1834
rect -782 1800 -748 1834
rect -690 1798 -656 1832
rect -572 1798 -538 1832
rect -386 1800 -352 1834
rect -270 1798 -236 1832
rect -178 1800 -144 1834
rect -14 1800 20 1834
rect 84 1798 118 1832
rect 242 1798 276 1832
rect 334 1798 368 1832
rect -1302 1188 -1268 1222
rect -1210 1188 -1176 1222
rect -1038 1188 -1004 1222
rect -936 1188 -902 1222
rect -784 1188 -750 1222
rect -690 1188 -656 1222
rect -564 1188 -530 1222
rect -386 1186 -352 1220
rect -270 1186 -236 1220
rect -178 1186 -144 1220
rect -14 1188 20 1222
rect 78 1186 112 1220
rect 242 1188 276 1222
rect 334 1186 368 1220
rect -478 1050 -444 1084
<< metal1 >>
rect -486 3008 -426 3012
rect -490 2956 -480 3008
rect -428 2956 -418 3008
rect -486 2824 -426 2956
rect -1410 2774 -578 2824
rect -588 2772 -578 2774
rect -526 2822 510 2824
rect -526 2774 514 2822
rect -526 2772 -516 2774
rect -1414 2728 -1360 2730
rect -878 2728 -868 2732
rect -1414 2680 -868 2728
rect -816 2728 -806 2732
rect -406 2728 -396 2730
rect -816 2680 -396 2728
rect -1414 2678 -396 2680
rect -344 2728 -334 2730
rect -106 2728 -96 2732
rect -344 2680 -96 2728
rect -44 2728 -34 2732
rect -44 2680 510 2728
rect -344 2678 510 2680
rect -1408 2582 508 2632
rect -700 2536 -690 2540
rect -1408 2488 -690 2536
rect -638 2536 -628 2540
rect -282 2536 -272 2538
rect -638 2488 -272 2536
rect -1408 2486 -272 2488
rect -220 2536 -210 2538
rect -220 2486 510 2536
rect 68 2440 78 2446
rect -1408 2438 78 2440
rect -1408 2390 -782 2438
rect -792 2386 -782 2390
rect -730 2394 78 2438
rect 130 2440 140 2446
rect 130 2394 508 2440
rect -730 2390 508 2394
rect -730 2386 -720 2390
rect -24 2344 -14 2348
rect -1408 2294 -950 2344
rect -960 2292 -950 2294
rect -898 2296 -14 2344
rect 38 2344 48 2348
rect 38 2296 508 2344
rect -898 2294 508 2296
rect -898 2292 -888 2294
rect -1050 2248 -1040 2250
rect -1408 2198 -1040 2248
rect -988 2248 -978 2250
rect -492 2248 -482 2250
rect -988 2198 -482 2248
rect -430 2248 -420 2250
rect -430 2198 508 2248
rect -1572 2082 -1332 2098
rect -1572 2030 -1510 2082
rect -1458 2030 -1332 2082
rect -1224 2034 -1214 2086
rect -1162 2034 -1152 2086
rect 230 2036 240 2088
rect 292 2036 302 2088
rect 392 2082 648 2102
rect -1572 2002 -1332 2030
rect 392 2030 524 2082
rect 576 2030 648 2082
rect 392 2006 648 2030
rect -496 1926 -486 1978
rect -434 1926 -424 1978
rect -1322 1788 -1312 1840
rect -1260 1788 -1250 1840
rect -1222 1788 -1212 1840
rect -1160 1788 -1150 1840
rect -1060 1794 -1050 1846
rect -998 1794 -988 1846
rect -960 1794 -950 1846
rect -898 1794 -888 1846
rect -804 1790 -794 1842
rect -742 1790 -732 1842
rect -704 1792 -694 1844
rect -642 1792 -632 1844
rect -590 1790 -580 1842
rect -528 1790 -518 1842
rect -404 1792 -394 1844
rect -342 1792 -332 1844
rect -290 1792 -280 1844
rect -228 1792 -218 1844
rect -190 1792 -180 1844
rect -128 1792 -118 1844
rect -32 1792 -22 1844
rect 30 1792 40 1844
rect 68 1792 78 1844
rect 130 1792 140 1844
rect 222 1790 232 1842
rect 284 1790 294 1842
rect 322 1790 332 1842
rect 384 1790 394 1842
rect -1316 1500 -1306 1552
rect -1254 1500 -1244 1552
rect -1224 1480 -1214 1532
rect -1162 1480 -1152 1532
rect 322 1506 332 1558
rect 384 1506 394 1558
rect -1326 1180 -1316 1232
rect -1264 1180 -1254 1232
rect -1224 1180 -1214 1232
rect -1162 1180 -1152 1232
rect -1058 1176 -1048 1228
rect -996 1176 -986 1228
rect -956 1178 -946 1230
rect -894 1178 -884 1230
rect -802 1180 -792 1232
rect -740 1180 -730 1232
rect -702 1180 -692 1232
rect -640 1180 -630 1232
rect -586 1178 -576 1230
rect -524 1178 -514 1230
rect -404 1178 -394 1230
rect -342 1178 -332 1230
rect -292 1180 -282 1232
rect -230 1180 -220 1232
rect -190 1180 -180 1232
rect -128 1180 -118 1232
rect -38 1178 -28 1230
rect 24 1178 34 1230
rect 66 1180 76 1232
rect 128 1180 138 1232
rect 216 1176 226 1228
rect 278 1176 288 1228
rect 322 1180 332 1232
rect 384 1180 394 1232
rect -496 1044 -486 1096
rect -434 1044 -424 1096
rect -1574 994 -1334 1016
rect 408 996 648 1014
rect -1574 942 -1510 994
rect -1458 942 -1334 994
rect -1320 944 -1310 996
rect -1258 944 -1248 996
rect 408 944 528 996
rect 580 944 648 996
rect -1574 920 -1334 942
rect 408 918 648 944
rect -1378 818 -574 822
rect -1378 770 -948 818
rect -958 766 -948 770
rect -896 770 -574 818
rect -522 770 420 822
rect -896 766 -886 770
rect -1380 718 426 724
rect -1380 666 -1130 718
rect -1078 712 426 718
rect -1078 666 -398 712
rect -1380 660 -398 666
rect -346 660 154 712
rect 206 660 426 712
rect -1376 606 420 614
rect -1376 554 -790 606
rect -738 554 -482 606
rect -430 554 420 606
rect -1376 550 420 554
rect -1378 492 422 504
rect -1378 440 -182 492
rect -130 440 -24 492
rect 28 440 422 492
rect -1380 382 424 394
rect -1380 330 -692 382
rect -640 330 -278 382
rect -226 330 424 382
rect -1382 282 238 284
rect -1382 230 78 282
rect 130 232 238 282
rect 290 232 424 284
rect 130 230 424 232
rect -1382 222 424 230
rect -1382 166 426 176
rect -1382 164 160 166
rect -1382 114 -1048 164
rect -1056 112 -1048 114
rect -996 114 160 164
rect 212 114 426 166
rect -996 112 -984 114
rect 384 68 426 70
rect -1382 58 426 68
rect -1382 6 -480 58
rect -428 6 332 58
rect 384 6 426 58
<< via1 >>
rect -480 2956 -428 3008
rect -578 2772 -526 2824
rect -868 2680 -816 2732
rect -396 2678 -344 2730
rect -96 2680 -44 2732
rect -690 2488 -638 2540
rect -272 2486 -220 2538
rect -782 2386 -730 2438
rect 78 2394 130 2446
rect -950 2292 -898 2344
rect -14 2296 38 2348
rect -1040 2198 -988 2250
rect -482 2198 -430 2250
rect -1510 2030 -1458 2082
rect -1214 2034 -1162 2086
rect 240 2036 292 2088
rect 524 2030 576 2082
rect -486 1970 -434 1978
rect -486 1936 -478 1970
rect -478 1936 -444 1970
rect -444 1936 -434 1970
rect -486 1926 -434 1936
rect -1312 1832 -1260 1840
rect -1312 1798 -1302 1832
rect -1302 1798 -1268 1832
rect -1268 1798 -1260 1832
rect -1312 1788 -1260 1798
rect -1212 1832 -1160 1840
rect -1212 1798 -1210 1832
rect -1210 1798 -1176 1832
rect -1176 1798 -1160 1832
rect -1212 1788 -1160 1798
rect -1050 1834 -998 1846
rect -1050 1800 -1038 1834
rect -1038 1800 -1004 1834
rect -1004 1800 -998 1834
rect -1050 1794 -998 1800
rect -950 1834 -898 1846
rect -950 1800 -946 1834
rect -946 1800 -912 1834
rect -912 1800 -898 1834
rect -950 1794 -898 1800
rect -794 1834 -742 1842
rect -794 1800 -782 1834
rect -782 1800 -748 1834
rect -748 1800 -742 1834
rect -794 1790 -742 1800
rect -694 1832 -642 1844
rect -694 1798 -690 1832
rect -690 1798 -656 1832
rect -656 1798 -642 1832
rect -694 1792 -642 1798
rect -580 1832 -528 1842
rect -580 1798 -572 1832
rect -572 1798 -538 1832
rect -538 1798 -528 1832
rect -580 1790 -528 1798
rect -394 1834 -342 1844
rect -394 1800 -386 1834
rect -386 1800 -352 1834
rect -352 1800 -342 1834
rect -394 1792 -342 1800
rect -280 1832 -228 1844
rect -280 1798 -270 1832
rect -270 1798 -236 1832
rect -236 1798 -228 1832
rect -280 1792 -228 1798
rect -180 1834 -128 1844
rect -180 1800 -178 1834
rect -178 1800 -144 1834
rect -144 1800 -128 1834
rect -180 1792 -128 1800
rect -22 1834 30 1844
rect -22 1800 -14 1834
rect -14 1800 20 1834
rect 20 1800 30 1834
rect -22 1792 30 1800
rect 78 1832 130 1844
rect 78 1798 84 1832
rect 84 1798 118 1832
rect 118 1798 130 1832
rect 78 1792 130 1798
rect 232 1832 284 1842
rect 232 1798 242 1832
rect 242 1798 276 1832
rect 276 1798 284 1832
rect 232 1790 284 1798
rect 332 1832 384 1842
rect 332 1798 334 1832
rect 334 1798 368 1832
rect 368 1798 384 1832
rect 332 1790 384 1798
rect -1306 1500 -1254 1552
rect -1214 1480 -1162 1532
rect 332 1506 384 1558
rect -1316 1222 -1264 1232
rect -1316 1188 -1302 1222
rect -1302 1188 -1268 1222
rect -1268 1188 -1264 1222
rect -1316 1180 -1264 1188
rect -1214 1222 -1162 1232
rect -1214 1188 -1210 1222
rect -1210 1188 -1176 1222
rect -1176 1188 -1162 1222
rect -1214 1180 -1162 1188
rect -1048 1222 -996 1228
rect -1048 1188 -1038 1222
rect -1038 1188 -1004 1222
rect -1004 1188 -996 1222
rect -1048 1176 -996 1188
rect -946 1222 -894 1230
rect -946 1188 -936 1222
rect -936 1188 -902 1222
rect -902 1188 -894 1222
rect -946 1178 -894 1188
rect -792 1222 -740 1232
rect -792 1188 -784 1222
rect -784 1188 -750 1222
rect -750 1188 -740 1222
rect -792 1180 -740 1188
rect -692 1222 -640 1232
rect -692 1188 -690 1222
rect -690 1188 -656 1222
rect -656 1188 -640 1222
rect -692 1180 -640 1188
rect -576 1222 -524 1230
rect -576 1188 -564 1222
rect -564 1188 -530 1222
rect -530 1188 -524 1222
rect -576 1178 -524 1188
rect -394 1220 -342 1230
rect -394 1186 -386 1220
rect -386 1186 -352 1220
rect -352 1186 -342 1220
rect -394 1178 -342 1186
rect -282 1220 -230 1232
rect -282 1186 -270 1220
rect -270 1186 -236 1220
rect -236 1186 -230 1220
rect -282 1180 -230 1186
rect -180 1220 -128 1232
rect -180 1186 -178 1220
rect -178 1186 -144 1220
rect -144 1186 -128 1220
rect -180 1180 -128 1186
rect -28 1222 24 1230
rect -28 1188 -14 1222
rect -14 1188 20 1222
rect 20 1188 24 1222
rect -28 1178 24 1188
rect 76 1220 128 1232
rect 76 1186 78 1220
rect 78 1186 112 1220
rect 112 1186 128 1220
rect 76 1180 128 1186
rect 226 1222 278 1228
rect 226 1188 242 1222
rect 242 1188 276 1222
rect 276 1188 278 1222
rect 226 1176 278 1188
rect 332 1220 384 1232
rect 332 1186 334 1220
rect 334 1186 368 1220
rect 368 1186 384 1220
rect 332 1180 384 1186
rect -486 1084 -434 1096
rect -486 1050 -478 1084
rect -478 1050 -444 1084
rect -444 1050 -434 1084
rect -486 1044 -434 1050
rect -1510 942 -1458 994
rect -1310 944 -1258 996
rect 528 944 580 996
rect -948 766 -896 818
rect -574 770 -522 822
rect -1130 666 -1078 718
rect -398 660 -346 712
rect 154 660 206 712
rect -790 554 -738 606
rect -482 554 -430 606
rect -182 440 -130 492
rect -24 440 28 492
rect -692 330 -640 382
rect -278 330 -226 382
rect 78 230 130 282
rect 238 232 290 284
rect -1048 112 -996 164
rect 160 114 212 166
rect -480 6 -428 58
rect 332 6 384 58
<< metal2 >>
rect -486 3012 -426 3022
rect -486 2942 -426 2952
rect -1134 2930 -1074 2940
rect -1410 2870 -1134 2904
rect 150 2932 210 2942
rect -1074 2872 150 2904
rect 210 2872 510 2904
rect -1074 2870 510 2872
rect -1134 2860 -1074 2870
rect -578 2824 -526 2834
rect -578 2762 -526 2772
rect -1510 2082 -1458 2092
rect -1510 994 -1458 2030
rect -1302 1850 -1256 2754
rect -1212 2096 -1166 2754
rect -1038 2260 -992 2754
rect -946 2354 -900 2754
rect -872 2738 -812 2748
rect -872 2668 -812 2678
rect -782 2448 -736 2754
rect -692 2550 -646 2754
rect -692 2540 -638 2550
rect -692 2488 -690 2540
rect -692 2478 -638 2488
rect -782 2438 -730 2448
rect -782 2376 -730 2386
rect -950 2344 -898 2354
rect -950 2282 -898 2292
rect -1040 2250 -988 2260
rect -1040 2188 -988 2198
rect -1214 2086 -1162 2096
rect -1214 2024 -1162 2034
rect -1312 1840 -1256 1850
rect -1260 1788 -1256 1840
rect -1312 1778 -1256 1788
rect -1302 1562 -1256 1778
rect -1212 1850 -1166 2024
rect -1038 1856 -992 2188
rect -946 1856 -900 2282
rect -1212 1840 -1160 1850
rect -1212 1778 -1160 1788
rect -1050 1846 -992 1856
rect -998 1794 -992 1846
rect -1050 1784 -992 1794
rect -950 1846 -898 1856
rect -782 1852 -736 2376
rect -692 1854 -646 2478
rect -950 1784 -898 1794
rect -794 1842 -736 1852
rect -742 1790 -736 1842
rect -1212 1576 -1166 1778
rect -1306 1552 -1254 1562
rect -1038 1558 -992 1784
rect -946 1558 -900 1784
rect -794 1780 -736 1790
rect -694 1844 -642 1854
rect -572 1852 -526 2762
rect -478 2260 -432 2754
rect -392 2740 -346 2754
rect -396 2730 -344 2740
rect -396 2668 -344 2678
rect -482 2250 -430 2260
rect -482 2188 -430 2198
rect -478 1988 -432 2188
rect -486 1978 -432 1988
rect -434 1926 -432 1978
rect -486 1916 -432 1926
rect -694 1782 -642 1792
rect -580 1842 -526 1852
rect -528 1790 -526 1842
rect -782 1558 -736 1780
rect -692 1558 -646 1782
rect -580 1780 -526 1790
rect -572 1558 -526 1780
rect -478 1558 -432 1916
rect -392 1854 -346 2668
rect -272 2548 -228 2754
rect -272 2538 -220 2548
rect -272 2476 -220 2486
rect -272 1854 -226 2476
rect -178 1854 -132 2870
rect 150 2862 210 2870
rect -102 2738 -42 2748
rect -102 2668 -42 2678
rect -14 2358 34 2754
rect 78 2456 124 2754
rect 78 2446 130 2456
rect 78 2384 130 2394
rect -14 2348 38 2358
rect -14 2286 38 2296
rect -14 1854 34 2286
rect -394 1844 -342 1854
rect -394 1782 -342 1792
rect -280 1844 -226 1854
rect -228 1792 -226 1844
rect -280 1782 -226 1792
rect -180 1844 -128 1854
rect -180 1782 -128 1792
rect -22 1844 34 1854
rect 30 1792 34 1844
rect -22 1782 34 1792
rect -392 1558 -346 1782
rect -272 1560 -226 1782
rect -178 1560 -132 1782
rect -14 1558 34 1782
rect 78 1854 124 2384
rect 242 2098 288 2754
rect 240 2088 292 2098
rect 240 2026 292 2036
rect 78 1844 130 1854
rect 242 1852 288 2026
rect 334 1852 380 2754
rect 524 2082 580 2092
rect 576 2030 580 2082
rect 524 2020 580 2030
rect 78 1782 130 1792
rect 232 1842 288 1852
rect 284 1790 288 1842
rect 78 1558 124 1782
rect 232 1780 288 1790
rect 332 1842 384 1852
rect 332 1780 384 1790
rect 242 1558 288 1780
rect 334 1568 380 1780
rect 332 1558 384 1568
rect -1306 1490 -1254 1500
rect -1214 1532 -1162 1542
rect 332 1496 384 1506
rect -1214 1470 -1162 1480
rect -1306 1242 -1260 1462
rect -1210 1242 -1164 1470
rect -1316 1232 -1260 1242
rect -1264 1180 -1260 1232
rect -1316 1170 -1260 1180
rect -1214 1232 -1162 1242
rect -1042 1238 -996 1462
rect -1214 1170 -1162 1180
rect -1048 1228 -996 1238
rect -1306 1006 -1260 1170
rect -1510 932 -1458 942
rect -1310 996 -1258 1006
rect -1310 934 -1258 944
rect -1306 146 -1260 934
rect -1210 146 -1164 1170
rect -1048 1166 -996 1176
rect -1134 722 -1074 732
rect -1134 652 -1074 662
rect -1042 180 -996 1166
rect -946 1240 -900 1462
rect -786 1242 -740 1462
rect -690 1242 -644 1462
rect -946 1230 -894 1240
rect -946 1168 -894 1178
rect -792 1232 -740 1242
rect -792 1170 -740 1180
rect -692 1232 -640 1242
rect -570 1240 -524 1464
rect -692 1170 -640 1180
rect -576 1230 -524 1240
rect -946 828 -900 1168
rect -786 836 -740 1170
rect -948 818 -896 828
rect -948 756 -896 766
rect -1050 170 -990 180
rect -946 146 -900 756
rect -790 616 -740 836
rect -790 606 -738 616
rect -790 544 -738 554
rect -790 540 -740 544
rect -790 146 -744 540
rect -690 392 -644 1170
rect -576 1168 -524 1178
rect -570 832 -524 1168
rect -478 1106 -432 1464
rect -486 1096 -432 1106
rect -434 1044 -432 1096
rect -486 1034 -432 1044
rect -574 822 -522 832
rect -574 760 -522 770
rect -692 382 -640 392
rect -692 320 -640 330
rect -690 146 -644 320
rect -570 146 -524 760
rect -478 616 -432 1034
rect -394 1240 -348 1464
rect -274 1242 -228 1462
rect -178 1242 -132 1462
rect -20 1276 26 1462
rect -394 1230 -342 1240
rect -394 1168 -342 1178
rect -282 1232 -228 1242
rect -230 1180 -228 1232
rect -282 1170 -228 1180
rect -180 1232 -128 1242
rect -22 1240 26 1276
rect 78 1242 124 1462
rect 240 1266 286 1462
rect -180 1170 -128 1180
rect -28 1230 26 1240
rect 24 1178 26 1230
rect -394 896 -348 1168
rect -396 722 -348 896
rect -398 712 -346 722
rect -398 650 -346 660
rect -482 606 -430 616
rect -482 544 -430 554
rect -478 146 -432 544
rect -396 146 -350 650
rect -274 392 -228 1170
rect -178 502 -132 1170
rect -28 1168 26 1178
rect 76 1232 128 1242
rect 240 1238 288 1266
rect 334 1242 382 1462
rect 76 1170 128 1180
rect 226 1228 288 1238
rect 278 1176 288 1228
rect -20 502 26 1168
rect 78 884 124 1170
rect 226 1166 288 1176
rect 332 1232 384 1242
rect 332 1170 384 1180
rect 78 750 126 884
rect 78 630 124 750
rect 152 716 212 726
rect 152 646 212 656
rect -182 492 -130 502
rect -182 430 -130 440
rect -24 492 28 502
rect -24 430 28 440
rect -278 382 -226 392
rect -278 320 -226 330
rect -274 146 -228 320
rect -178 146 -132 430
rect -20 146 26 430
rect 78 292 126 630
rect 240 294 288 1166
rect 78 282 130 292
rect 78 220 130 230
rect 238 284 290 294
rect 238 222 290 232
rect 78 148 126 220
rect 240 208 288 222
rect 80 146 126 148
rect 154 170 214 180
rect -1050 100 -990 110
rect 242 146 288 208
rect 154 100 214 110
rect -486 62 -426 72
rect 334 68 382 1170
rect 528 996 580 2020
rect 528 934 580 944
rect -486 -8 -426 2
rect 332 58 384 68
rect 332 -4 384 6
<< via2 >>
rect -486 3008 -426 3012
rect -486 2956 -480 3008
rect -480 2956 -428 3008
rect -428 2956 -426 3008
rect -486 2952 -426 2956
rect -1134 2870 -1074 2930
rect 150 2872 210 2932
rect -872 2732 -812 2738
rect -872 2680 -868 2732
rect -868 2680 -816 2732
rect -816 2680 -812 2732
rect -872 2678 -812 2680
rect -102 2732 -42 2738
rect -102 2680 -96 2732
rect -96 2680 -44 2732
rect -44 2680 -42 2732
rect -102 2678 -42 2680
rect -1134 718 -1074 722
rect -1134 666 -1130 718
rect -1130 666 -1078 718
rect -1078 666 -1074 718
rect -1134 662 -1074 666
rect -1050 164 -990 170
rect -1050 112 -1048 164
rect -1048 112 -996 164
rect -996 112 -990 164
rect 152 712 212 716
rect 152 660 154 712
rect 154 660 206 712
rect 206 660 212 712
rect 152 656 212 660
rect 154 166 214 170
rect -1050 110 -990 112
rect 154 114 160 166
rect 160 114 212 166
rect 212 114 214 166
rect 154 110 214 114
rect -486 58 -426 62
rect -486 6 -480 58
rect -480 6 -428 58
rect -428 6 -426 58
rect -486 2 -426 6
<< metal3 >>
rect -496 3012 -416 3018
rect -496 2952 -486 3012
rect -426 2952 -416 3012
rect -1144 2930 -1064 2940
rect -1144 2870 -1134 2930
rect -1074 2870 -1064 2930
rect -1144 722 -1064 2870
rect -1144 662 -1134 722
rect -1074 662 -1064 722
rect -1144 656 -1064 662
rect -912 2744 -832 2940
rect -912 2738 -802 2744
rect -912 2678 -872 2738
rect -812 2678 -802 2738
rect -912 2673 -802 2678
rect -1060 174 -980 175
rect -912 174 -832 2673
rect -1060 170 -832 174
rect -1060 110 -1050 170
rect -990 110 -832 170
rect -1060 100 -832 110
rect -496 62 -416 2952
rect -82 2748 -2 2954
rect 142 2937 222 2940
rect 140 2932 222 2937
rect 140 2872 150 2932
rect 210 2872 222 2932
rect 140 2867 222 2872
rect -112 2738 0 2748
rect -112 2678 -102 2738
rect -42 2678 0 2738
rect -112 2670 0 2678
rect -82 174 -2 2670
rect 142 716 222 2867
rect 142 656 152 716
rect 212 656 222 716
rect 142 646 222 656
rect 144 174 224 175
rect -82 170 224 174
rect -82 110 154 170
rect 214 110 224 170
rect -82 105 224 110
rect -82 100 162 105
rect -82 94 -2 100
rect -496 2 -486 62
rect -426 2 -416 62
rect -496 -12 -416 2
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 -854 0 1 966
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1676037725
transform 1 0 -342 0 1 966
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1676037725
transform 1 0 -86 0 1 966
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1676037725
transform 1 0 170 0 1 966
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1676037725
transform 1 0 170 0 -1 2054
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1676037725
transform 1 0 -1110 0 1 966
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1676037725
transform -1 0 -1098 0 -1 2054
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1676037725
transform 1 0 -1110 0 -1 2054
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1676037725
transform 1 0 -854 0 -1 2054
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1676037725
transform 1 0 -342 0 -1 2054
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_11
timestamp 1676037725
transform 1 0 -86 0 -1 2054
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_12
timestamp 1676037725
transform 1 0 -1374 0 1 966
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 -598 0 -1 2054
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_2
timestamp 1676037725
transform 1 0 -598 0 1 966
box -38 -48 314 592
<< labels >>
rlabel metal1 474 2216 474 2216 1 net1
rlabel metal1 464 2302 464 2302 1 net2
rlabel metal1 466 2404 466 2404 1 net3
rlabel metal2 460 2882 460 2882 1 net5
rlabel metal1 -1364 790 -1364 790 1 net4
rlabel metal1 -1366 572 -1366 572 1 net6
rlabel metal1 -1366 344 -1366 344 1 net7
rlabel metal1 -1366 464 -1366 464 1 net8
rlabel metal1 -1366 12 -1366 12 1 net9
flabel metal1 -1382 222 -1382 222 1 FreeSans 160 0 0 0 do_clk2_1v8
port 3 n
flabel metal2 550 1118 550 1118 1 FreeSans 160 0 0 0 VSS_CG
port 1 n
flabel locali -1604 1484 -1604 1484 1 FreeSans 160 0 0 0 VDD_CG
port 4 n
flabel metal1 -1408 2486 -1408 2486 1 FreeSans 160 0 0 0 do_clk1_1v8
port 2 n
flabel metal1 -1382 114 -1370 120 1 FreeSans 160 0 0 0 di_clk_1v8
port 0 n
<< end >>
