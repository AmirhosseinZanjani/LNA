magic
tech sky130A
magscale 1 2
timestamp 1710847391
<< nwell >>
rect -12515 -1219 12515 1219
<< pmos >>
rect -12319 -1000 -10319 1000
rect -10261 -1000 -8261 1000
rect -8203 -1000 -6203 1000
rect -6145 -1000 -4145 1000
rect -4087 -1000 -2087 1000
rect -2029 -1000 -29 1000
rect 29 -1000 2029 1000
rect 2087 -1000 4087 1000
rect 4145 -1000 6145 1000
rect 6203 -1000 8203 1000
rect 8261 -1000 10261 1000
rect 10319 -1000 12319 1000
<< pdiff >>
rect -12377 988 -12319 1000
rect -12377 -988 -12365 988
rect -12331 -988 -12319 988
rect -12377 -1000 -12319 -988
rect -10319 988 -10261 1000
rect -10319 -988 -10307 988
rect -10273 -988 -10261 988
rect -10319 -1000 -10261 -988
rect -8261 988 -8203 1000
rect -8261 -988 -8249 988
rect -8215 -988 -8203 988
rect -8261 -1000 -8203 -988
rect -6203 988 -6145 1000
rect -6203 -988 -6191 988
rect -6157 -988 -6145 988
rect -6203 -1000 -6145 -988
rect -4145 988 -4087 1000
rect -4145 -988 -4133 988
rect -4099 -988 -4087 988
rect -4145 -1000 -4087 -988
rect -2087 988 -2029 1000
rect -2087 -988 -2075 988
rect -2041 -988 -2029 988
rect -2087 -1000 -2029 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 2029 988 2087 1000
rect 2029 -988 2041 988
rect 2075 -988 2087 988
rect 2029 -1000 2087 -988
rect 4087 988 4145 1000
rect 4087 -988 4099 988
rect 4133 -988 4145 988
rect 4087 -1000 4145 -988
rect 6145 988 6203 1000
rect 6145 -988 6157 988
rect 6191 -988 6203 988
rect 6145 -1000 6203 -988
rect 8203 988 8261 1000
rect 8203 -988 8215 988
rect 8249 -988 8261 988
rect 8203 -1000 8261 -988
rect 10261 988 10319 1000
rect 10261 -988 10273 988
rect 10307 -988 10319 988
rect 10261 -1000 10319 -988
rect 12319 988 12377 1000
rect 12319 -988 12331 988
rect 12365 -988 12377 988
rect 12319 -1000 12377 -988
<< pdiffc >>
rect -12365 -988 -12331 988
rect -10307 -988 -10273 988
rect -8249 -988 -8215 988
rect -6191 -988 -6157 988
rect -4133 -988 -4099 988
rect -2075 -988 -2041 988
rect -17 -988 17 988
rect 2041 -988 2075 988
rect 4099 -988 4133 988
rect 6157 -988 6191 988
rect 8215 -988 8249 988
rect 10273 -988 10307 988
rect 12331 -988 12365 988
<< nsubdiff >>
rect -12479 1149 -12383 1183
rect 12383 1149 12479 1183
rect -12479 1087 -12445 1149
rect 12445 1087 12479 1149
rect -12479 -1149 -12445 -1087
rect 12445 -1149 12479 -1087
rect -12479 -1183 -12383 -1149
rect 12383 -1183 12479 -1149
<< nsubdiffcont >>
rect -12383 1149 12383 1183
rect -12479 -1087 -12445 1087
rect 12445 -1087 12479 1087
rect -12383 -1183 12383 -1149
<< poly >>
rect -12319 1081 -10319 1097
rect -12319 1047 -12303 1081
rect -10335 1047 -10319 1081
rect -12319 1000 -10319 1047
rect -10261 1081 -8261 1097
rect -10261 1047 -10245 1081
rect -8277 1047 -8261 1081
rect -10261 1000 -8261 1047
rect -8203 1081 -6203 1097
rect -8203 1047 -8187 1081
rect -6219 1047 -6203 1081
rect -8203 1000 -6203 1047
rect -6145 1081 -4145 1097
rect -6145 1047 -6129 1081
rect -4161 1047 -4145 1081
rect -6145 1000 -4145 1047
rect -4087 1081 -2087 1097
rect -4087 1047 -4071 1081
rect -2103 1047 -2087 1081
rect -4087 1000 -2087 1047
rect -2029 1081 -29 1097
rect -2029 1047 -2013 1081
rect -45 1047 -29 1081
rect -2029 1000 -29 1047
rect 29 1081 2029 1097
rect 29 1047 45 1081
rect 2013 1047 2029 1081
rect 29 1000 2029 1047
rect 2087 1081 4087 1097
rect 2087 1047 2103 1081
rect 4071 1047 4087 1081
rect 2087 1000 4087 1047
rect 4145 1081 6145 1097
rect 4145 1047 4161 1081
rect 6129 1047 6145 1081
rect 4145 1000 6145 1047
rect 6203 1081 8203 1097
rect 6203 1047 6219 1081
rect 8187 1047 8203 1081
rect 6203 1000 8203 1047
rect 8261 1081 10261 1097
rect 8261 1047 8277 1081
rect 10245 1047 10261 1081
rect 8261 1000 10261 1047
rect 10319 1081 12319 1097
rect 10319 1047 10335 1081
rect 12303 1047 12319 1081
rect 10319 1000 12319 1047
rect -12319 -1047 -10319 -1000
rect -12319 -1081 -12303 -1047
rect -10335 -1081 -10319 -1047
rect -12319 -1097 -10319 -1081
rect -10261 -1047 -8261 -1000
rect -10261 -1081 -10245 -1047
rect -8277 -1081 -8261 -1047
rect -10261 -1097 -8261 -1081
rect -8203 -1047 -6203 -1000
rect -8203 -1081 -8187 -1047
rect -6219 -1081 -6203 -1047
rect -8203 -1097 -6203 -1081
rect -6145 -1047 -4145 -1000
rect -6145 -1081 -6129 -1047
rect -4161 -1081 -4145 -1047
rect -6145 -1097 -4145 -1081
rect -4087 -1047 -2087 -1000
rect -4087 -1081 -4071 -1047
rect -2103 -1081 -2087 -1047
rect -4087 -1097 -2087 -1081
rect -2029 -1047 -29 -1000
rect -2029 -1081 -2013 -1047
rect -45 -1081 -29 -1047
rect -2029 -1097 -29 -1081
rect 29 -1047 2029 -1000
rect 29 -1081 45 -1047
rect 2013 -1081 2029 -1047
rect 29 -1097 2029 -1081
rect 2087 -1047 4087 -1000
rect 2087 -1081 2103 -1047
rect 4071 -1081 4087 -1047
rect 2087 -1097 4087 -1081
rect 4145 -1047 6145 -1000
rect 4145 -1081 4161 -1047
rect 6129 -1081 6145 -1047
rect 4145 -1097 6145 -1081
rect 6203 -1047 8203 -1000
rect 6203 -1081 6219 -1047
rect 8187 -1081 8203 -1047
rect 6203 -1097 8203 -1081
rect 8261 -1047 10261 -1000
rect 8261 -1081 8277 -1047
rect 10245 -1081 10261 -1047
rect 8261 -1097 10261 -1081
rect 10319 -1047 12319 -1000
rect 10319 -1081 10335 -1047
rect 12303 -1081 12319 -1047
rect 10319 -1097 12319 -1081
<< polycont >>
rect -12303 1047 -10335 1081
rect -10245 1047 -8277 1081
rect -8187 1047 -6219 1081
rect -6129 1047 -4161 1081
rect -4071 1047 -2103 1081
rect -2013 1047 -45 1081
rect 45 1047 2013 1081
rect 2103 1047 4071 1081
rect 4161 1047 6129 1081
rect 6219 1047 8187 1081
rect 8277 1047 10245 1081
rect 10335 1047 12303 1081
rect -12303 -1081 -10335 -1047
rect -10245 -1081 -8277 -1047
rect -8187 -1081 -6219 -1047
rect -6129 -1081 -4161 -1047
rect -4071 -1081 -2103 -1047
rect -2013 -1081 -45 -1047
rect 45 -1081 2013 -1047
rect 2103 -1081 4071 -1047
rect 4161 -1081 6129 -1047
rect 6219 -1081 8187 -1047
rect 8277 -1081 10245 -1047
rect 10335 -1081 12303 -1047
<< locali >>
rect -12479 1149 -12383 1183
rect 12383 1149 12479 1183
rect -12479 1087 -12445 1149
rect 12445 1087 12479 1149
rect -12319 1047 -12303 1081
rect -10335 1047 -10319 1081
rect -10261 1047 -10245 1081
rect -8277 1047 -8261 1081
rect -8203 1047 -8187 1081
rect -6219 1047 -6203 1081
rect -6145 1047 -6129 1081
rect -4161 1047 -4145 1081
rect -4087 1047 -4071 1081
rect -2103 1047 -2087 1081
rect -2029 1047 -2013 1081
rect -45 1047 -29 1081
rect 29 1047 45 1081
rect 2013 1047 2029 1081
rect 2087 1047 2103 1081
rect 4071 1047 4087 1081
rect 4145 1047 4161 1081
rect 6129 1047 6145 1081
rect 6203 1047 6219 1081
rect 8187 1047 8203 1081
rect 8261 1047 8277 1081
rect 10245 1047 10261 1081
rect 10319 1047 10335 1081
rect 12303 1047 12319 1081
rect -12365 988 -12331 1004
rect -12365 -1004 -12331 -988
rect -10307 988 -10273 1004
rect -10307 -1004 -10273 -988
rect -8249 988 -8215 1004
rect -8249 -1004 -8215 -988
rect -6191 988 -6157 1004
rect -6191 -1004 -6157 -988
rect -4133 988 -4099 1004
rect -4133 -1004 -4099 -988
rect -2075 988 -2041 1004
rect -2075 -1004 -2041 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 2041 988 2075 1004
rect 2041 -1004 2075 -988
rect 4099 988 4133 1004
rect 4099 -1004 4133 -988
rect 6157 988 6191 1004
rect 6157 -1004 6191 -988
rect 8215 988 8249 1004
rect 8215 -1004 8249 -988
rect 10273 988 10307 1004
rect 10273 -1004 10307 -988
rect 12331 988 12365 1004
rect 12331 -1004 12365 -988
rect -12319 -1081 -12303 -1047
rect -10335 -1081 -10319 -1047
rect -10261 -1081 -10245 -1047
rect -8277 -1081 -8261 -1047
rect -8203 -1081 -8187 -1047
rect -6219 -1081 -6203 -1047
rect -6145 -1081 -6129 -1047
rect -4161 -1081 -4145 -1047
rect -4087 -1081 -4071 -1047
rect -2103 -1081 -2087 -1047
rect -2029 -1081 -2013 -1047
rect -45 -1081 -29 -1047
rect 29 -1081 45 -1047
rect 2013 -1081 2029 -1047
rect 2087 -1081 2103 -1047
rect 4071 -1081 4087 -1047
rect 4145 -1081 4161 -1047
rect 6129 -1081 6145 -1047
rect 6203 -1081 6219 -1047
rect 8187 -1081 8203 -1047
rect 8261 -1081 8277 -1047
rect 10245 -1081 10261 -1047
rect 10319 -1081 10335 -1047
rect 12303 -1081 12319 -1047
rect -12479 -1149 -12445 -1087
rect 12445 -1149 12479 -1087
rect -12479 -1183 -12383 -1149
rect 12383 -1183 12479 -1149
<< viali >>
rect -12303 1047 -10335 1081
rect -10245 1047 -8277 1081
rect -8187 1047 -6219 1081
rect -6129 1047 -4161 1081
rect -4071 1047 -2103 1081
rect -2013 1047 -45 1081
rect 45 1047 2013 1081
rect 2103 1047 4071 1081
rect 4161 1047 6129 1081
rect 6219 1047 8187 1081
rect 8277 1047 10245 1081
rect 10335 1047 12303 1081
rect -12365 -988 -12331 988
rect -10307 -988 -10273 988
rect -8249 -988 -8215 988
rect -6191 -988 -6157 988
rect -4133 -988 -4099 988
rect -2075 -988 -2041 988
rect -17 -988 17 988
rect 2041 -988 2075 988
rect 4099 -988 4133 988
rect 6157 -988 6191 988
rect 8215 -988 8249 988
rect 10273 -988 10307 988
rect 12331 -988 12365 988
rect -12303 -1081 -10335 -1047
rect -10245 -1081 -8277 -1047
rect -8187 -1081 -6219 -1047
rect -6129 -1081 -4161 -1047
rect -4071 -1081 -2103 -1047
rect -2013 -1081 -45 -1047
rect 45 -1081 2013 -1047
rect 2103 -1081 4071 -1047
rect 4161 -1081 6129 -1047
rect 6219 -1081 8187 -1047
rect 8277 -1081 10245 -1047
rect 10335 -1081 12303 -1047
<< metal1 >>
rect -12315 1081 -10323 1087
rect -12315 1047 -12303 1081
rect -10335 1047 -10323 1081
rect -12315 1041 -10323 1047
rect -10257 1081 -8265 1087
rect -10257 1047 -10245 1081
rect -8277 1047 -8265 1081
rect -10257 1041 -8265 1047
rect -8199 1081 -6207 1087
rect -8199 1047 -8187 1081
rect -6219 1047 -6207 1081
rect -8199 1041 -6207 1047
rect -6141 1081 -4149 1087
rect -6141 1047 -6129 1081
rect -4161 1047 -4149 1081
rect -6141 1041 -4149 1047
rect -4083 1081 -2091 1087
rect -4083 1047 -4071 1081
rect -2103 1047 -2091 1081
rect -4083 1041 -2091 1047
rect -2025 1081 -33 1087
rect -2025 1047 -2013 1081
rect -45 1047 -33 1081
rect -2025 1041 -33 1047
rect 33 1081 2025 1087
rect 33 1047 45 1081
rect 2013 1047 2025 1081
rect 33 1041 2025 1047
rect 2091 1081 4083 1087
rect 2091 1047 2103 1081
rect 4071 1047 4083 1081
rect 2091 1041 4083 1047
rect 4149 1081 6141 1087
rect 4149 1047 4161 1081
rect 6129 1047 6141 1081
rect 4149 1041 6141 1047
rect 6207 1081 8199 1087
rect 6207 1047 6219 1081
rect 8187 1047 8199 1081
rect 6207 1041 8199 1047
rect 8265 1081 10257 1087
rect 8265 1047 8277 1081
rect 10245 1047 10257 1081
rect 8265 1041 10257 1047
rect 10323 1081 12315 1087
rect 10323 1047 10335 1081
rect 12303 1047 12315 1081
rect 10323 1041 12315 1047
rect -12371 988 -12325 1000
rect -12371 -988 -12365 988
rect -12331 -988 -12325 988
rect -12371 -1000 -12325 -988
rect -10313 988 -10267 1000
rect -10313 -988 -10307 988
rect -10273 -988 -10267 988
rect -10313 -1000 -10267 -988
rect -8255 988 -8209 1000
rect -8255 -988 -8249 988
rect -8215 -988 -8209 988
rect -8255 -1000 -8209 -988
rect -6197 988 -6151 1000
rect -6197 -988 -6191 988
rect -6157 -988 -6151 988
rect -6197 -1000 -6151 -988
rect -4139 988 -4093 1000
rect -4139 -988 -4133 988
rect -4099 -988 -4093 988
rect -4139 -1000 -4093 -988
rect -2081 988 -2035 1000
rect -2081 -988 -2075 988
rect -2041 -988 -2035 988
rect -2081 -1000 -2035 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 2035 988 2081 1000
rect 2035 -988 2041 988
rect 2075 -988 2081 988
rect 2035 -1000 2081 -988
rect 4093 988 4139 1000
rect 4093 -988 4099 988
rect 4133 -988 4139 988
rect 4093 -1000 4139 -988
rect 6151 988 6197 1000
rect 6151 -988 6157 988
rect 6191 -988 6197 988
rect 6151 -1000 6197 -988
rect 8209 988 8255 1000
rect 8209 -988 8215 988
rect 8249 -988 8255 988
rect 8209 -1000 8255 -988
rect 10267 988 10313 1000
rect 10267 -988 10273 988
rect 10307 -988 10313 988
rect 10267 -1000 10313 -988
rect 12325 988 12371 1000
rect 12325 -988 12331 988
rect 12365 -988 12371 988
rect 12325 -1000 12371 -988
rect -12315 -1047 -10323 -1041
rect -12315 -1081 -12303 -1047
rect -10335 -1081 -10323 -1047
rect -12315 -1087 -10323 -1081
rect -10257 -1047 -8265 -1041
rect -10257 -1081 -10245 -1047
rect -8277 -1081 -8265 -1047
rect -10257 -1087 -8265 -1081
rect -8199 -1047 -6207 -1041
rect -8199 -1081 -8187 -1047
rect -6219 -1081 -6207 -1047
rect -8199 -1087 -6207 -1081
rect -6141 -1047 -4149 -1041
rect -6141 -1081 -6129 -1047
rect -4161 -1081 -4149 -1047
rect -6141 -1087 -4149 -1081
rect -4083 -1047 -2091 -1041
rect -4083 -1081 -4071 -1047
rect -2103 -1081 -2091 -1047
rect -4083 -1087 -2091 -1081
rect -2025 -1047 -33 -1041
rect -2025 -1081 -2013 -1047
rect -45 -1081 -33 -1047
rect -2025 -1087 -33 -1081
rect 33 -1047 2025 -1041
rect 33 -1081 45 -1047
rect 2013 -1081 2025 -1047
rect 33 -1087 2025 -1081
rect 2091 -1047 4083 -1041
rect 2091 -1081 2103 -1047
rect 4071 -1081 4083 -1047
rect 2091 -1087 4083 -1081
rect 4149 -1047 6141 -1041
rect 4149 -1081 4161 -1047
rect 6129 -1081 6141 -1047
rect 4149 -1087 6141 -1081
rect 6207 -1047 8199 -1041
rect 6207 -1081 6219 -1047
rect 8187 -1081 8199 -1047
rect 6207 -1087 8199 -1081
rect 8265 -1047 10257 -1041
rect 8265 -1081 8277 -1047
rect 10245 -1081 10257 -1047
rect 8265 -1087 10257 -1081
rect 10323 -1047 12315 -1041
rect 10323 -1081 10335 -1047
rect 12303 -1081 12315 -1047
rect 10323 -1087 12315 -1081
<< properties >>
string FIXED_BBOX -12462 -1166 12462 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 10 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
