magic
tech sky130A
magscale 1 2
timestamp 1710866800
<< viali >>
rect 24889 3480 24941 3532
rect 88 1361 140 1413
rect 1116 1361 1168 1413
rect 23754 1361 23806 1413
rect 24784 1361 24836 1413
<< metal1 >>
rect 1106 3590 1116 3642
rect 1168 3590 1178 3642
rect 3164 3590 3174 3642
rect 3226 3590 3236 3642
rect 5226 3592 5236 3644
rect 5288 3592 5298 3644
rect 7280 3588 7290 3640
rect 7342 3588 7352 3640
rect 9338 3590 9348 3642
rect 9400 3590 9410 3642
rect 11396 3590 11406 3642
rect 11458 3590 11468 3642
rect 13454 3590 13464 3642
rect 13516 3590 13526 3642
rect 15512 3590 15522 3642
rect 15574 3590 15584 3642
rect 17570 3590 17580 3642
rect 17632 3590 17642 3642
rect 19628 3590 19638 3642
rect 19690 3590 19700 3642
rect 21686 3590 21696 3642
rect 21748 3590 21758 3642
rect 23744 3590 23754 3642
rect 23806 3590 23816 3642
rect 24877 3532 24953 3538
rect 78 3480 88 3532
rect 140 3480 150 3532
rect 2136 3480 2146 3532
rect 2198 3480 2208 3532
rect 4194 3480 4204 3532
rect 4256 3480 4266 3532
rect 6252 3480 6262 3532
rect 6314 3480 6324 3532
rect 8310 3480 8320 3532
rect 8372 3480 8382 3532
rect 10368 3480 10378 3532
rect 10430 3480 10440 3532
rect 12426 3480 12436 3532
rect 12488 3480 12498 3532
rect 14484 3480 14494 3532
rect 14546 3480 14556 3532
rect 16540 3480 16550 3532
rect 16602 3480 16612 3532
rect 18602 3480 18612 3532
rect 18664 3480 18674 3532
rect 20658 3480 20668 3532
rect 20720 3480 20730 3532
rect 22716 3480 22726 3532
rect 22778 3480 22788 3532
rect 24774 3480 24784 3532
rect 24836 3480 24846 3532
rect 24877 3480 24889 3532
rect 24941 3480 24953 3532
rect 24877 3474 24953 3480
rect 78 1556 88 1608
rect 140 1556 150 1608
rect 2136 1556 2146 1608
rect 2198 1556 2208 1608
rect 4194 1556 4204 1608
rect 4256 1556 4266 1608
rect 6252 1556 6262 1608
rect 6314 1556 6324 1608
rect 8310 1556 8320 1608
rect 8372 1556 8382 1608
rect 10368 1556 10378 1608
rect 10430 1556 10440 1608
rect 12426 1556 12436 1608
rect 12488 1556 12498 1608
rect 14484 1556 14494 1608
rect 14546 1556 14556 1608
rect 16540 1556 16550 1608
rect 16602 1556 16612 1608
rect 18600 1556 18610 1608
rect 18662 1556 18672 1608
rect 20658 1556 20668 1608
rect 20720 1556 20730 1608
rect 22716 1556 22726 1608
rect 22778 1556 22788 1608
rect 24774 1556 24784 1608
rect 24836 1556 24846 1608
rect 24879 1556 24889 1608
rect 24941 1556 24951 1608
rect 1106 1462 1116 1514
rect 1168 1462 1178 1514
rect 3164 1462 3174 1514
rect 3226 1462 3236 1514
rect 5226 1460 5236 1512
rect 5288 1460 5298 1512
rect 7280 1460 7290 1512
rect 7342 1460 7352 1512
rect 9338 1462 9348 1514
rect 9400 1462 9410 1514
rect 11396 1462 11406 1514
rect 11458 1462 11468 1514
rect 13454 1462 13464 1514
rect 13516 1462 13526 1514
rect 15512 1462 15522 1514
rect 15574 1462 15584 1514
rect 17570 1462 17580 1514
rect 17632 1462 17642 1514
rect 19628 1462 19638 1514
rect 19690 1462 19700 1514
rect 21686 1462 21696 1514
rect 21748 1462 21758 1514
rect 23744 1462 23754 1514
rect 23806 1462 23816 1514
rect 76 1413 152 1419
rect 76 1361 88 1413
rect 140 1361 152 1413
rect 76 1355 152 1361
rect 1104 1413 1180 1419
rect 1104 1361 1116 1413
rect 1168 1361 1180 1413
rect 1104 1355 1180 1361
rect 23742 1413 23818 1419
rect 23742 1361 23754 1413
rect 23806 1361 23818 1413
rect 23742 1355 23818 1361
rect 24772 1413 24848 1419
rect 24772 1361 24784 1413
rect 24836 1361 24848 1413
rect 24772 1355 24848 1361
<< via1 >>
rect 1116 3590 1168 3642
rect 3174 3590 3226 3642
rect 5236 3592 5288 3644
rect 7290 3588 7342 3640
rect 9348 3590 9400 3642
rect 11406 3590 11458 3642
rect 13464 3590 13516 3642
rect 15522 3590 15574 3642
rect 17580 3590 17632 3642
rect 19638 3590 19690 3642
rect 21696 3590 21748 3642
rect 23754 3590 23806 3642
rect 88 3480 140 3532
rect 2146 3480 2198 3532
rect 4204 3480 4256 3532
rect 6262 3480 6314 3532
rect 8320 3480 8372 3532
rect 10378 3480 10430 3532
rect 12436 3480 12488 3532
rect 14494 3480 14546 3532
rect 16550 3480 16602 3532
rect 18612 3480 18664 3532
rect 20668 3480 20720 3532
rect 22726 3480 22778 3532
rect 24784 3480 24836 3532
rect 24889 3480 24941 3532
rect 88 1556 140 1608
rect 2146 1556 2198 1608
rect 4204 1556 4256 1608
rect 6262 1556 6314 1608
rect 8320 1556 8372 1608
rect 10378 1556 10430 1608
rect 12436 1556 12488 1608
rect 14494 1556 14546 1608
rect 16550 1556 16602 1608
rect 18610 1556 18662 1608
rect 20668 1556 20720 1608
rect 22726 1556 22778 1608
rect 24784 1556 24836 1608
rect 24889 1556 24941 1608
rect 1116 1462 1168 1514
rect 3174 1462 3226 1514
rect 5236 1460 5288 1512
rect 7290 1460 7342 1512
rect 9348 1462 9400 1514
rect 11406 1462 11458 1514
rect 13464 1462 13516 1514
rect 15522 1462 15574 1514
rect 17580 1462 17632 1514
rect 19638 1462 19690 1514
rect 21696 1462 21748 1514
rect 23754 1462 23806 1514
rect 88 1361 140 1413
rect 1116 1361 1168 1413
rect 23754 1361 23806 1413
rect 24784 1361 24836 1413
<< metal2 >>
rect 88 3532 140 3727
rect -17 3480 88 3532
rect 88 1608 140 3480
rect -17 1556 88 1608
rect 88 1413 140 1556
rect 88 620 140 1361
rect 1116 3642 1168 4174
rect 3174 3898 3226 4174
rect 5236 4022 5288 4174
rect 5234 4012 5292 4022
rect 5234 3946 5292 3956
rect 3170 3888 3228 3898
rect 3170 3822 3228 3832
rect 1116 1514 1168 3590
rect 3174 3642 3226 3822
rect 1116 1413 1168 1462
rect 1116 1351 1168 1361
rect 2146 3532 2198 3542
rect 2146 1608 2198 3480
rect 2146 1266 2198 1556
rect 3174 1514 3226 3590
rect 5236 3644 5288 3946
rect 7290 3898 7342 4174
rect 9348 4022 9400 4174
rect 9346 4012 9404 4022
rect 9346 3946 9404 3956
rect 7286 3888 7344 3898
rect 7286 3822 7344 3832
rect 3174 1452 3226 1462
rect 4204 3532 4256 3542
rect 4204 1608 4256 3480
rect 2144 1256 2202 1266
rect 2144 1190 2202 1200
rect 2146 620 2198 1190
rect 4204 1140 4256 1556
rect 5236 1512 5288 3592
rect 7290 3640 7342 3822
rect 5236 1450 5288 1460
rect 6262 3532 6314 3542
rect 6262 1608 6314 3480
rect 4200 1130 4258 1140
rect 4200 1064 4258 1074
rect 4204 620 4256 1064
rect 6262 1016 6314 1556
rect 7290 1512 7342 3588
rect 9348 3642 9400 3946
rect 11406 3898 11458 4174
rect 13464 4022 13516 4174
rect 13460 4012 13518 4022
rect 13460 3946 13518 3956
rect 11404 3888 11462 3898
rect 11404 3822 11462 3832
rect 7290 1450 7342 1460
rect 8320 3532 8372 3542
rect 8320 1608 8372 3480
rect 8320 1140 8372 1556
rect 9348 1514 9400 3590
rect 11406 3642 11458 3822
rect 9348 1452 9400 1462
rect 10378 3532 10430 3542
rect 10378 1608 10430 3480
rect 10378 1266 10430 1556
rect 11406 1514 11458 3590
rect 13464 3642 13516 3946
rect 15522 3898 15574 4174
rect 17580 4022 17632 4174
rect 17576 4012 17634 4022
rect 17576 3946 17634 3956
rect 15520 3888 15578 3898
rect 15520 3822 15578 3832
rect 11406 1452 11458 1462
rect 12436 3532 12488 3542
rect 12436 1608 12488 3480
rect 10376 1256 10434 1266
rect 10376 1190 10434 1200
rect 8316 1130 8374 1140
rect 8316 1064 8374 1074
rect 6260 1006 6318 1016
rect 6260 940 6318 950
rect 6262 620 6314 940
rect 8320 620 8372 1064
rect 10378 620 10430 1190
rect 12436 1140 12488 1556
rect 13464 1514 13516 3590
rect 15522 3642 15574 3822
rect 13464 1452 13516 1462
rect 14494 3532 14546 3542
rect 14494 1608 14546 3480
rect 12432 1130 12490 1140
rect 12432 1064 12490 1074
rect 12436 620 12488 1064
rect 14494 1016 14546 1556
rect 15522 1514 15574 3590
rect 17580 3642 17632 3946
rect 19638 3898 19690 4174
rect 21696 4022 21748 4174
rect 21694 4012 21752 4022
rect 21694 3946 21752 3956
rect 19634 3888 19692 3898
rect 19634 3822 19692 3832
rect 15522 1452 15574 1462
rect 16550 3532 16602 3542
rect 16550 1608 16602 3480
rect 16550 1140 16602 1556
rect 17580 1514 17632 3590
rect 19638 3642 19690 3822
rect 18612 3532 18664 3542
rect 18612 3470 18664 3480
rect 18612 2298 18662 3470
rect 17580 1452 17632 1462
rect 18610 1608 18662 2298
rect 18610 1266 18662 1556
rect 19638 1514 19690 3590
rect 21696 3642 21748 3946
rect 19638 1452 19690 1462
rect 20668 3532 20720 3542
rect 20668 1608 20720 3480
rect 18606 1256 18664 1266
rect 18606 1190 18664 1200
rect 16546 1130 16604 1140
rect 16546 1064 16604 1074
rect 14492 1006 14550 1016
rect 14492 940 14550 950
rect 14494 620 14546 940
rect 16550 620 16602 1064
rect 18610 620 18662 1190
rect 20668 1140 20720 1556
rect 21696 1514 21748 3590
rect 23754 3642 23806 4174
rect 21696 1452 21748 1462
rect 22726 3532 22778 3542
rect 22726 1608 22778 3480
rect 20664 1130 20722 1140
rect 20664 1064 20722 1074
rect 20668 620 20720 1064
rect 22726 1016 22778 1556
rect 23754 1514 23806 3590
rect 23754 1413 23806 1462
rect 23754 1351 23806 1361
rect 24784 3532 24836 3727
rect 24889 3532 24941 3542
rect 24836 3480 24889 3532
rect 24784 1608 24836 3480
rect 24889 3470 24941 3480
rect 24889 1608 24941 1618
rect 24836 1556 24889 1608
rect 24784 1413 24836 1556
rect 24889 1546 24941 1556
rect 22724 1006 22782 1016
rect 22724 940 22782 950
rect 22726 620 22778 940
rect 24784 620 24836 1361
<< via2 >>
rect 5234 3956 5292 4012
rect 3170 3832 3228 3888
rect 9346 3956 9404 4012
rect 7286 3832 7344 3888
rect 2144 1200 2202 1256
rect 4200 1074 4258 1130
rect 13460 3956 13518 4012
rect 11404 3832 11462 3888
rect 17576 3956 17634 4012
rect 15520 3832 15578 3888
rect 10376 1200 10434 1256
rect 8316 1074 8374 1130
rect 6260 950 6318 1006
rect 12432 1074 12490 1130
rect 21694 3956 21752 4012
rect 19634 3832 19692 3888
rect 18606 1200 18664 1256
rect 16546 1074 16604 1130
rect 14492 950 14550 1006
rect 20664 1074 20722 1130
rect 22724 950 22782 1006
<< metal3 >>
rect -54 4078 25702 4138
rect 5224 4014 5302 4017
rect 9336 4014 9414 4017
rect 13450 4014 13528 4017
rect 17566 4014 17644 4017
rect 21684 4014 21762 4017
rect -54 4012 25702 4014
rect -54 3956 5234 4012
rect 5292 3956 9346 4012
rect 9404 3956 13460 4012
rect 13518 3956 17576 4012
rect 17634 3956 21694 4012
rect 21752 3956 25702 4012
rect -54 3954 25702 3956
rect 5224 3951 5302 3954
rect 9336 3951 9414 3954
rect 13450 3951 13528 3954
rect 17566 3951 17644 3954
rect 21684 3951 21762 3954
rect 3160 3890 3238 3893
rect 7276 3890 7354 3893
rect 11394 3890 11472 3893
rect 15510 3890 15588 3893
rect 19624 3890 19702 3893
rect -54 3888 25702 3890
rect -54 3832 3170 3888
rect 3228 3832 7286 3888
rect 7344 3832 11404 3888
rect 11462 3832 15520 3888
rect 15578 3832 19634 3888
rect 19692 3832 25702 3888
rect -54 3830 25702 3832
rect 3160 3827 3238 3830
rect 7276 3827 7354 3830
rect 11394 3827 11472 3830
rect 15510 3827 15588 3830
rect 19624 3827 19702 3830
rect 2134 1258 2212 1261
rect 10366 1258 10444 1261
rect 18596 1258 18674 1261
rect -126 1256 25630 1258
rect -126 1200 2144 1256
rect 2202 1200 10376 1256
rect 10434 1200 18606 1256
rect 18664 1200 25630 1256
rect -126 1198 25630 1200
rect -126 1196 3300 1198
rect 2134 1195 2212 1196
rect 10366 1195 10444 1198
rect 18596 1195 18674 1198
rect 4190 1132 4268 1135
rect 8306 1132 8384 1135
rect 12422 1132 12500 1135
rect 16536 1132 16614 1135
rect 20654 1132 20732 1135
rect -126 1130 25630 1132
rect -126 1074 4200 1130
rect 4258 1074 8316 1130
rect 8374 1074 12432 1130
rect 12490 1074 16546 1130
rect 16604 1074 20664 1130
rect 20722 1074 25630 1130
rect -126 1072 25630 1074
rect 4190 1069 4268 1072
rect 8306 1069 8384 1072
rect 12422 1069 12500 1072
rect 16536 1069 16614 1072
rect 20654 1069 20732 1072
rect 6250 1008 6328 1011
rect 14482 1008 14560 1011
rect 22714 1008 22792 1011
rect -126 1006 25630 1008
rect -126 950 6260 1006
rect 6318 950 14492 1006
rect 14550 950 22724 1006
rect 22782 950 25630 1006
rect -126 948 25630 950
rect 6250 945 6328 948
rect 14482 945 14560 948
rect 22714 945 22792 948
use sky130_fd_pr__pfet_01v8_X3BJMD  sky130_fd_pr__pfet_01v8_X3BJMD_0
timestamp 1710847391
transform 1 0 12462 0 1 2544
box -12515 -1219 12515 1219
<< end >>
