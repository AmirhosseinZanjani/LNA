magic
tech sky130A
magscale 1 2
timestamp 1710869429
<< viali >>
rect -437698 1962556 -437646 1962608
<< metal1 >>
rect -460346 1964889 -460336 1964941
rect -460284 1964889 -460274 1964941
rect -437708 1964889 -437698 1964941
rect -437646 1964889 -437636 1964941
rect -460347 1964787 -460337 1964839
rect -460285 1964787 -460275 1964839
rect -458288 1964786 -458278 1964838
rect -458226 1964786 -458216 1964838
rect -456229 1964787 -456219 1964839
rect -456167 1964787 -456157 1964839
rect -454172 1964787 -454162 1964839
rect -454110 1964787 -454100 1964839
rect -452116 1964787 -452106 1964839
rect -452054 1964787 -452044 1964839
rect -450056 1964786 -450046 1964838
rect -449994 1964786 -449984 1964838
rect -447998 1964786 -447988 1964838
rect -447936 1964786 -447926 1964838
rect -445939 1964785 -445929 1964837
rect -445877 1964785 -445867 1964837
rect -443883 1964786 -443873 1964838
rect -443821 1964786 -443811 1964838
rect -441824 1964785 -441814 1964837
rect -441762 1964785 -441752 1964837
rect -439766 1964787 -439756 1964839
rect -439704 1964787 -439694 1964839
rect -437708 1964786 -437698 1964838
rect -437646 1964786 -437636 1964838
rect -461375 1964676 -461365 1964728
rect -461313 1964676 -461303 1964728
rect -459317 1964676 -459307 1964728
rect -459255 1964676 -459245 1964728
rect -457258 1964676 -457248 1964728
rect -457196 1964676 -457186 1964728
rect -455201 1964676 -455191 1964728
rect -455139 1964676 -455129 1964728
rect -453143 1964676 -453133 1964728
rect -453081 1964676 -453071 1964728
rect -451084 1964676 -451074 1964728
rect -451022 1964676 -451012 1964728
rect -449027 1964676 -449017 1964728
rect -448965 1964676 -448955 1964728
rect -446969 1964676 -446959 1964728
rect -446907 1964676 -446897 1964728
rect -444911 1964676 -444901 1964728
rect -444849 1964676 -444839 1964728
rect -442853 1964677 -442843 1964729
rect -442791 1964677 -442781 1964729
rect -440795 1964677 -440785 1964729
rect -440733 1964677 -440723 1964729
rect -438738 1964676 -438728 1964728
rect -438676 1964676 -438666 1964728
rect -436679 1964676 -436669 1964728
rect -436617 1964676 -436607 1964728
rect -461375 1962752 -461365 1962804
rect -461313 1962752 -461303 1962804
rect -459317 1962752 -459307 1962804
rect -459255 1962752 -459245 1962804
rect -457258 1962752 -457248 1962804
rect -457196 1962752 -457186 1962804
rect -455201 1962752 -455191 1962804
rect -455139 1962752 -455129 1962804
rect -453143 1962752 -453133 1962804
rect -453081 1962752 -453071 1962804
rect -451085 1962752 -451075 1962804
rect -451023 1962752 -451013 1962804
rect -449027 1962752 -449017 1962804
rect -448965 1962752 -448955 1962804
rect -446969 1962752 -446959 1962804
rect -446907 1962752 -446897 1962804
rect -444910 1962752 -444900 1962804
rect -444848 1962752 -444838 1962804
rect -442852 1962752 -442842 1962804
rect -442790 1962752 -442780 1962804
rect -440796 1962752 -440786 1962804
rect -440734 1962752 -440724 1962804
rect -438736 1962752 -438726 1962804
rect -438674 1962752 -438664 1962804
rect -436679 1962752 -436669 1962804
rect -436617 1962752 -436607 1962804
rect -460346 1962659 -460336 1962711
rect -460284 1962659 -460274 1962711
rect -458287 1962659 -458277 1962711
rect -458225 1962659 -458215 1962711
rect -456229 1962659 -456219 1962711
rect -456167 1962659 -456157 1962711
rect -454172 1962659 -454162 1962711
rect -454110 1962659 -454100 1962711
rect -452114 1962659 -452104 1962711
rect -452052 1962659 -452042 1962711
rect -450056 1962659 -450046 1962711
rect -449994 1962659 -449984 1962711
rect -447998 1962659 -447988 1962711
rect -447936 1962659 -447926 1962711
rect -445940 1962659 -445930 1962711
rect -445878 1962659 -445868 1962711
rect -443882 1962659 -443872 1962711
rect -443820 1962659 -443810 1962711
rect -441824 1962659 -441814 1962711
rect -441762 1962659 -441752 1962711
rect -439766 1962660 -439756 1962712
rect -439704 1962660 -439694 1962712
rect -437708 1962659 -437698 1962711
rect -437646 1962659 -437636 1962711
rect -460346 1962557 -460336 1962609
rect -460284 1962557 -460274 1962609
rect -437710 1962608 -437634 1962614
rect -437710 1962556 -437698 1962608
rect -437646 1962556 -437634 1962608
rect -437710 1962550 -437634 1962556
<< via1 >>
rect -460336 1964889 -460284 1964941
rect -437698 1964889 -437646 1964941
rect -460337 1964787 -460285 1964839
rect -458278 1964786 -458226 1964838
rect -456219 1964787 -456167 1964839
rect -454162 1964787 -454110 1964839
rect -452106 1964787 -452054 1964839
rect -450046 1964786 -449994 1964838
rect -447988 1964786 -447936 1964838
rect -445929 1964785 -445877 1964837
rect -443873 1964786 -443821 1964838
rect -441814 1964785 -441762 1964837
rect -439756 1964787 -439704 1964839
rect -437698 1964786 -437646 1964838
rect -461365 1964676 -461313 1964728
rect -459307 1964676 -459255 1964728
rect -457248 1964676 -457196 1964728
rect -455191 1964676 -455139 1964728
rect -453133 1964676 -453081 1964728
rect -451074 1964676 -451022 1964728
rect -449017 1964676 -448965 1964728
rect -446959 1964676 -446907 1964728
rect -444901 1964676 -444849 1964728
rect -442843 1964677 -442791 1964729
rect -440785 1964677 -440733 1964729
rect -438728 1964676 -438676 1964728
rect -436669 1964676 -436617 1964728
rect -461365 1962752 -461313 1962804
rect -459307 1962752 -459255 1962804
rect -457248 1962752 -457196 1962804
rect -455191 1962752 -455139 1962804
rect -453133 1962752 -453081 1962804
rect -451075 1962752 -451023 1962804
rect -449017 1962752 -448965 1962804
rect -446959 1962752 -446907 1962804
rect -444900 1962752 -444848 1962804
rect -442842 1962752 -442790 1962804
rect -440786 1962752 -440734 1962804
rect -438726 1962752 -438674 1962804
rect -436669 1962752 -436617 1962804
rect -460336 1962659 -460284 1962711
rect -458277 1962659 -458225 1962711
rect -456219 1962659 -456167 1962711
rect -454162 1962659 -454110 1962711
rect -452104 1962659 -452052 1962711
rect -450046 1962659 -449994 1962711
rect -447988 1962659 -447936 1962711
rect -445930 1962659 -445878 1962711
rect -443872 1962659 -443820 1962711
rect -441814 1962659 -441762 1962711
rect -439756 1962660 -439704 1962712
rect -437698 1962659 -437646 1962711
rect -460336 1962557 -460284 1962609
rect -437698 1962556 -437646 1962608
<< metal2 >>
rect -460336 1964941 -460284 1965497
rect -458277 1965092 -458225 1965497
rect -458280 1965082 -458224 1965092
rect -456219 1965091 -456167 1965497
rect -458280 1965016 -458224 1965026
rect -456223 1965081 -456167 1965091
rect -454162 1965090 -454110 1965497
rect -452104 1965092 -452052 1965497
rect -450046 1965092 -449994 1965497
rect -447988 1965093 -447936 1965497
rect -460336 1964849 -460284 1964889
rect -460337 1964839 -460284 1964849
rect -458277 1964848 -458225 1965016
rect -456223 1965015 -456167 1965025
rect -460285 1964787 -460284 1964839
rect -460337 1964777 -460284 1964787
rect -461469 1964738 -461322 1964744
rect -461469 1964728 -461313 1964738
rect -461469 1964676 -461365 1964728
rect -461365 1962805 -461313 1964676
rect -461470 1962804 -461311 1962805
rect -461470 1962803 -461365 1962804
rect -461471 1962752 -461365 1962803
rect -461313 1962752 -461311 1962804
rect -461471 1962737 -461311 1962752
rect -461471 1962735 -461313 1962737
rect -461365 1961871 -461313 1962735
rect -460336 1962711 -460284 1964777
rect -458278 1964838 -458225 1964848
rect -458226 1964786 -458225 1964838
rect -458278 1964776 -458225 1964786
rect -459298 1964738 -459264 1964744
rect -460336 1962609 -460284 1962659
rect -460336 1962547 -460284 1962557
rect -459307 1964728 -459255 1964738
rect -459307 1962804 -459255 1964676
rect -459307 1962496 -459255 1962752
rect -458277 1962711 -458225 1964776
rect -456219 1964839 -456167 1965015
rect -454166 1965080 -454110 1965090
rect -454166 1965014 -454110 1965024
rect -452107 1965082 -452051 1965092
rect -452107 1965016 -452051 1965026
rect -450049 1965082 -449993 1965092
rect -450049 1965016 -449993 1965026
rect -447991 1965083 -447935 1965093
rect -445930 1965091 -445878 1965497
rect -443872 1965092 -443821 1965497
rect -441814 1965092 -441762 1965497
rect -439756 1965093 -439704 1965497
rect -447991 1965017 -447935 1965027
rect -445933 1965081 -445877 1965091
rect -458277 1962649 -458225 1962659
rect -457248 1964728 -457196 1964738
rect -457248 1962804 -457196 1964676
rect -459308 1962146 -459255 1962496
rect -457248 1962366 -457196 1962752
rect -456219 1962711 -456167 1964787
rect -454162 1964839 -454110 1965014
rect -452104 1964849 -452052 1965016
rect -456219 1962649 -456167 1962659
rect -455191 1964728 -455139 1964744
rect -455191 1964666 -455139 1964676
rect -455191 1962814 -455140 1964666
rect -455191 1962804 -455139 1962814
rect -459308 1962090 -459256 1962146
rect -459309 1962080 -459253 1962090
rect -459309 1962014 -459253 1962024
rect -459308 1961871 -459256 1962014
rect -457248 1961964 -457195 1962366
rect -455191 1962233 -455139 1962752
rect -454162 1962711 -454110 1964787
rect -452106 1964839 -452052 1964849
rect -452054 1964787 -452052 1964839
rect -452106 1964777 -452052 1964787
rect -453133 1964728 -453081 1964738
rect -453133 1962814 -453081 1964676
rect -454162 1962649 -454110 1962659
rect -453136 1962804 -453081 1962814
rect -453136 1962752 -453133 1962804
rect -453136 1962742 -453081 1962752
rect -453136 1962372 -453084 1962742
rect -452104 1962711 -452052 1964777
rect -450046 1964838 -449994 1965016
rect -451074 1964735 -451022 1964738
rect -452104 1962649 -452052 1962659
rect -451075 1964728 -451022 1964735
rect -451075 1964676 -451074 1964728
rect -451075 1962804 -451022 1964676
rect -451023 1962752 -451022 1962804
rect -453137 1962250 -453083 1962372
rect -455192 1962090 -455139 1962233
rect -453139 1962199 -453083 1962250
rect -453138 1962146 -453083 1962199
rect -455194 1962080 -455138 1962090
rect -455194 1962014 -455138 1962024
rect -457251 1961954 -457195 1961964
rect -457251 1961888 -457195 1961898
rect -457248 1961077 -457195 1961888
rect -455192 1961871 -455140 1962014
rect -453138 1961964 -453084 1962146
rect -451075 1962090 -451022 1962752
rect -450046 1962711 -449994 1964786
rect -447988 1964838 -447936 1965017
rect -445933 1965015 -445877 1965025
rect -443876 1965082 -443820 1965092
rect -443876 1965016 -443820 1965026
rect -441818 1965082 -441762 1965092
rect -441818 1965016 -441762 1965026
rect -439760 1965083 -439704 1965093
rect -439760 1965017 -439704 1965027
rect -450046 1962649 -449994 1962659
rect -449017 1964728 -448965 1964738
rect -449017 1962804 -448965 1964676
rect -448965 1962752 -448964 1962753
rect -449017 1962378 -448964 1962752
rect -447988 1962711 -447936 1964786
rect -445930 1964847 -445878 1965015
rect -443872 1964848 -443821 1965016
rect -445930 1964837 -445877 1964847
rect -445930 1964785 -445929 1964837
rect -445930 1964775 -445877 1964785
rect -443873 1964838 -443821 1964848
rect -443873 1964776 -443821 1964786
rect -446959 1964728 -446907 1964738
rect -446959 1964666 -446907 1964676
rect -446959 1962804 -446907 1962814
rect -447988 1962649 -447936 1962659
rect -446963 1962752 -446959 1962753
rect -446963 1962742 -446907 1962752
rect -449017 1962146 -448963 1962378
rect -446963 1962247 -446910 1962742
rect -445930 1962711 -445878 1964775
rect -444901 1964728 -444849 1964738
rect -444901 1964666 -444849 1964676
rect -444900 1962804 -444848 1962814
rect -444900 1962746 -444848 1962752
rect -445930 1962649 -445878 1962659
rect -444904 1962742 -444848 1962746
rect -451078 1962080 -451022 1962090
rect -451078 1962014 -451022 1962024
rect -453141 1961954 -453084 1961964
rect -453141 1961888 -453085 1961898
rect -453138 1961077 -453085 1961888
rect -451075 1961871 -451022 1962014
rect -449016 1961965 -448963 1962146
rect -446964 1962090 -446910 1962247
rect -446966 1962080 -446910 1962090
rect -446966 1962014 -446910 1962024
rect -449018 1961955 -448962 1961965
rect -449018 1961889 -448962 1961899
rect -449016 1961077 -448963 1961889
rect -446964 1961871 -446910 1962014
rect -444904 1961965 -444851 1962742
rect -443872 1962721 -443821 1964776
rect -441814 1964837 -441762 1965016
rect -442843 1964729 -442791 1964739
rect -442843 1964667 -442791 1964677
rect -442842 1962804 -442790 1962814
rect -442845 1962752 -442842 1962753
rect -442845 1962742 -442790 1962752
rect -443872 1962711 -443820 1962721
rect -443872 1962649 -443820 1962659
rect -442845 1962203 -442792 1962742
rect -441814 1962711 -441762 1964785
rect -439756 1964839 -439704 1965017
rect -440785 1964729 -440733 1964739
rect -440785 1964667 -440733 1964677
rect -440786 1962804 -440734 1962814
rect -441814 1962649 -441762 1962659
rect -440790 1962752 -440786 1962753
rect -440790 1962742 -440734 1962752
rect -442846 1962090 -442792 1962203
rect -442848 1962080 -442792 1962090
rect -442848 1962014 -442792 1962024
rect -444907 1961955 -444851 1961965
rect -444907 1961889 -444851 1961899
rect -444904 1961077 -444851 1961889
rect -442846 1961871 -442792 1962014
rect -440790 1962361 -440737 1962742
rect -439756 1962712 -439704 1964787
rect -437698 1965140 -437645 1965497
rect -437698 1964941 -437643 1965140
rect -437646 1964889 -437645 1964941
rect -437698 1964838 -437645 1964889
rect -437646 1964786 -437645 1964838
rect -438728 1964728 -438676 1964738
rect -438728 1964666 -438676 1964676
rect -438726 1962804 -438674 1962814
rect -439756 1962650 -439704 1962660
rect -438728 1962752 -438726 1962753
rect -438728 1962742 -438674 1962752
rect -440790 1961965 -440736 1962361
rect -438728 1962090 -438675 1962742
rect -437698 1962711 -437645 1964786
rect -436669 1964728 -436512 1964744
rect -436617 1964676 -436512 1964728
rect -436669 1964666 -436617 1964676
rect -436669 1962804 -436617 1962814
rect -437646 1962659 -437645 1962711
rect -437698 1962608 -437645 1962659
rect -437646 1962556 -437645 1962608
rect -436672 1962752 -436669 1962753
rect -436617 1962752 -436512 1962804
rect -436672 1962736 -436512 1962752
rect -437698 1962546 -437646 1962556
rect -436672 1962228 -436619 1962736
rect -438733 1962080 -438675 1962090
rect -438677 1962024 -438675 1962080
rect -438733 1962014 -438675 1962024
rect -440792 1961955 -440736 1961965
rect -440792 1961889 -440736 1961899
rect -440790 1961077 -440736 1961889
rect -438728 1961871 -438675 1962014
rect -436673 1961871 -436618 1962228
<< via2 >>
rect -458280 1965026 -458224 1965082
rect -456223 1965025 -456167 1965081
rect -454166 1965024 -454110 1965080
rect -452107 1965026 -452051 1965082
rect -450049 1965026 -449993 1965082
rect -447991 1965027 -447935 1965083
rect -445933 1965025 -445877 1965081
rect -459309 1962024 -459253 1962080
rect -455194 1962024 -455138 1962080
rect -457251 1961898 -457195 1961954
rect -443876 1965026 -443820 1965082
rect -441818 1965026 -441762 1965082
rect -439760 1965027 -439704 1965083
rect -451078 1962024 -451022 1962080
rect -453141 1961898 -453085 1961954
rect -446966 1962024 -446910 1962080
rect -449018 1961899 -448962 1961955
rect -442848 1962024 -442792 1962080
rect -444907 1961899 -444851 1961955
rect -438733 1962024 -438677 1962080
rect -440792 1961899 -440736 1961955
<< metal3 >>
rect -461366 1965396 -436613 1965457
rect -461366 1965271 -436613 1965332
rect -461366 1965148 -436613 1965211
rect -461540 1965086 -460183 1965087
rect -458290 1965086 -458214 1965087
rect -452117 1965086 -452041 1965087
rect -450059 1965086 -449983 1965087
rect -448001 1965086 -447925 1965088
rect -443886 1965086 -443810 1965087
rect -441828 1965086 -441752 1965087
rect -439770 1965086 -437543 1965088
rect -461540 1965083 -436441 1965086
rect -461540 1965082 -447991 1965083
rect -461540 1965026 -458280 1965082
rect -458224 1965081 -452107 1965082
rect -458224 1965026 -456223 1965081
rect -461540 1965025 -456223 1965026
rect -456167 1965080 -452107 1965081
rect -456167 1965025 -454166 1965080
rect -461540 1965024 -454166 1965025
rect -454110 1965026 -452107 1965080
rect -452051 1965026 -450049 1965082
rect -449993 1965027 -447991 1965082
rect -447935 1965082 -439760 1965083
rect -447935 1965081 -443876 1965082
rect -447935 1965027 -445933 1965081
rect -449993 1965026 -445933 1965027
rect -454110 1965025 -445933 1965026
rect -445877 1965026 -443876 1965081
rect -443820 1965026 -441818 1965082
rect -441762 1965027 -439760 1965082
rect -439704 1965027 -436441 1965083
rect -441762 1965026 -436441 1965027
rect -445877 1965025 -436441 1965026
rect -454110 1965024 -436441 1965025
rect -461540 1965023 -436441 1965024
rect -458290 1965021 -458214 1965023
rect -456233 1965020 -456157 1965023
rect -454176 1965019 -454100 1965023
rect -452117 1965021 -452041 1965023
rect -450059 1965021 -449983 1965023
rect -448001 1965022 -447925 1965023
rect -445943 1965020 -445867 1965023
rect -443886 1965021 -443810 1965023
rect -441828 1965021 -441752 1965023
rect -439770 1965022 -439694 1965023
rect -461371 1962459 -438543 1962462
rect -461371 1962396 -436613 1962459
rect -461369 1962334 -444741 1962336
rect -461369 1962333 -440679 1962334
rect -461369 1962270 -436613 1962333
rect -461369 1962146 -436613 1962209
rect -461540 1962082 -459772 1962083
rect -459319 1962082 -459243 1962085
rect -455204 1962082 -455128 1962085
rect -451088 1962082 -451012 1962085
rect -446976 1962082 -446900 1962085
rect -442858 1962082 -442782 1962085
rect -438743 1962082 -438667 1962085
rect -461540 1962080 -436441 1962082
rect -461540 1962024 -459309 1962080
rect -459253 1962024 -455194 1962080
rect -455138 1962024 -451078 1962080
rect -451022 1962024 -446966 1962080
rect -446910 1962024 -442848 1962080
rect -442792 1962024 -438733 1962080
rect -438677 1962024 -436441 1962080
rect -461540 1962022 -436441 1962024
rect -461369 1962021 -436441 1962022
rect -459319 1962019 -459243 1962021
rect -455204 1962019 -455128 1962021
rect -451088 1962019 -451012 1962021
rect -446976 1962019 -446900 1962021
rect -442858 1962019 -442782 1962021
rect -438743 1962019 -438667 1962021
rect -457261 1961957 -457185 1961959
rect -453151 1961957 -453075 1961959
rect -449028 1961957 -448952 1961960
rect -444917 1961957 -444841 1961960
rect -440802 1961957 -440726 1961960
rect -461540 1961955 -436441 1961957
rect -461540 1961954 -449018 1961955
rect -461540 1961898 -457251 1961954
rect -457195 1961898 -453141 1961954
rect -453085 1961899 -449018 1961954
rect -448962 1961899 -444907 1961955
rect -444851 1961899 -440792 1961955
rect -440736 1961899 -436441 1961955
rect -453085 1961898 -436441 1961899
rect -461540 1961896 -436441 1961898
rect -457261 1961893 -457185 1961896
rect -453151 1961893 -453075 1961896
rect -449028 1961894 -448952 1961896
rect -444917 1961894 -444841 1961896
rect -440802 1961894 -440726 1961896
use sky130_fd_pr__pfet_01v8_X3BJMD  sky130_fd_pr__pfet_01v8_X3BJMD_0
timestamp 1710847391
transform 1 0 -448991 0 1 1963740
box -12515 -1219 12515 1219
<< end >>
